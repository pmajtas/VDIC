/******************************************************************************
 * (C) Copyright 2022 AGH UST All Rights Reserved
 ******************************************************************************
 * MODULE NAME: vdic_dut_2022
 * VERSION:     1.1
 * DATE:        03-11-2022
 *
 * ABSTRACT:   DUT module for VDIC 2022 labs.
 *              The DUT is RPN calculator type. The arguments are sent first,
 *              than the operator/command.
 *******************************************************************************
 * INPUTS
 *    clk      - posedge active clock, always running
 *    rst_n    - synchronous reset active low
 *    din      - serial data input
 *    enable_n - chip enable, active low;

 * OUTPUTS
 *    dout       - serial data output
 *    dout_valid - valid flag for serial data output, active high
 *
 *******************************************************************************

 The clock is always active.
 The DUT operates on the posedge of the clock.
 The DUT receives the data when enable_n is active.

 --------------------------------------------------------------------------------
 --- Input data
 --------------------------------------------------------------------------------

 The input data is send serially in WORDs.

 The WORD is always 10 bit long. MSB is sent first.
 The WORD sent to the DUT is either DATA type or CONTROL type.

 DATA = 0bbbbbbbbp
 where:
 - b = 0 or 1, PAYLOAD bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 CONTROL = 1bbbbbbbbp
 where:
 - b = 0 or 1, COMMAND bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 The COMMAND can be:
 00000000 - CMD_NOP, do nothing, remove the data (reset data stack)
 00000001 - CMD_AND, logic AND of the last two arguments
 00000010 - CMD_OR, logic OR of the arguments
 00000011 - CMD_XOR, logic XOR of the arguments
 00010000 - CMD_ADD, add the arguments
 00100000 - CMD_SUB, subtract other arguments from the first one

 --------------------------------------------------------------------------------
 --- Output data
 --------------------------------------------------------------------------------

 The DUT responds to each CONTROL word, sending 3 WORDS:
 STATUS, DATA, DATA

 STATUS = 1bbbbbbbbp
 where bbbbbbbb is one of:

 00000000 - S_NO_ERROR - data correctly processed
 00000001 - S_MISSING_DATA - missing input data
 00000010 - S_DATA_STACK_OVERFLOW - maximum number of arguments exceeded
 00000100 - S_OUTPUT_FIFO_OVERFLOW - result dropped not possible to process
 00100000 - S_DATA_PARITY_ERROR - input data or command parity error
 01000000 - S_COMMAND_PARITY_ERROR - input data or command parity error
 10000000 - S_INVALID_COMMAND - unknown command detected

 DATA is defined as in the input.
 PAYLOAD of the DATA is 00000000 if the data was NOT processed correctly.

 *******************************************************************************
 * IMPLEMENTATION STATUS
 *******************************************************************************
 *  <Feature>                        <Is implemented>
 *    command CMD_NOP                   YES
 *    command CMD_AND                   YES
 *    command CMD_OR                    YES
 *    command CMD_XOR                   YES
 *    command CMD_ADD                   YES
 *    command CMD_SUB                   YES
 *    status S_NO_ERROR                 YES
 *    status S_MISSING_DATA              NO
 *    status S_DATA_STACK_OVERFLOW       NO
 *    status S_OUTPUT_FIFO_OVERFLOW      NO
 *    status S_DATA_PARITY_ERROR         NO
 *    status S_COMMAND_PARITY_ERROR      NO
 *    status S_INVALID_COMMAND          YES
 *******************************************************************************
 */

// Generated by Cadence Genus(TM) Synthesis Solution 19.15-s090_1
// Generated on: Nov  3 2022 14:33:56 CET (Nov  3 2022 13:33:56 UTC)

// Verification Directory ./LEC 

module vdic_dut_2022(clk, rst_n, enable_n, din, dout, dout_valid);
  input clk, rst_n, enable_n, din;
  output dout, dout_valid;
  wire clk, rst_n, enable_n, din;
  wire dout, dout_valid;
  wire [7:0] \data_stack_mem[0] ;
  wire [7:0] \data_stack_mem[1] ;
  wire [7:0] \data_stack_mem[2] ;
  wire [7:0] \data_stack_mem[3] ;
  wire [7:0] \data_stack_mem[4] ;
  wire [7:0] \data_stack_mem[5] ;
  wire [7:0] \data_stack_mem[6] ;
  wire [7:0] \data_stack_mem[7] ;
  wire [7:0] \data_stack_mem[8] ;
  wire [3:0] data_stack_pointer;
  wire [3:0] sh_bit_cnt;
  wire [9:0] sh_reg_in;
  wire [4:0] sh_reg_out_bit_counter;
  wire [2:0] out_fifo_write_pointer;
  wire [2:0] out_fifo_read_pointer;
  wire [9:0] \out_fifo[6][0] ;
  wire [9:0] \out_fifo[3][0] ;
  wire [9:0] \out_fifo[7][0] ;
  wire [9:0] \out_fifo[0][0] ;
  wire [9:0] \out_fifo[4][0] ;
  wire [9:0] \out_fifo[2][0] ;
  wire [9:0] \out_fifo[4][1] ;
  wire [9:0] \out_fifo[5][2] ;
  wire [9:0] \out_fifo[2][2] ;
  wire [9:0] \out_fifo[1][2] ;
  wire [9:0] \out_fifo[6][2] ;
  wire [9:0] \out_fifo[3][2] ;
  wire [9:0] \out_fifo[7][2] ;
  wire [9:0] \out_fifo[0][2] ;
  wire [9:0] \out_fifo[4][2] ;
  wire [9:0] \out_fifo[1][1] ;
  wire [9:0] \out_fifo[7][1] ;
  wire [9:0] \out_fifo[0][1] ;
  wire [9:0] \out_fifo[5][0] ;
  wire [9:0] \out_fifo[3][1] ;
  wire [9:0] \out_fifo[6][1] ;
  wire [9:0] \out_fifo[1][0] ;
  wire [9:0] \out_fifo[2][1] ;
  wire [9:0] \out_fifo[5][1] ;
  wire [29:0] sh_reg_out;
  wire n_13813, n_13814, n_13815, n_13816, n_13823, n_13824, n_13825,
       n_13826;
  wire n_13827, n_13828, n_13829, n_13830, n_13831, n_13832, n_13833,
       n_13834;
  wire n_13835, n_13836, n_13837, n_13838, n_13839, n_13840, n_13841,
       n_13842;
  wire n_13843, n_13844, n_13845, n_13846, n_13847, n_13850, n_13851,
       n_13853;
  wire n_13854, n_13855, n_13856, n_13857, n_13858, n_13859, n_13860,
       n_13861;
  wire n_13862, n_13863, n_13864, n_13865, n_13866, n_13867, n_13868,
       n_13869;
  wire n_13870, n_13871, n_13872, n_13873, n_13874, n_13875, n_13876,
       n_13877;
  wire n_13878, n_13879, n_13880, n_13881, n_13882, n_13883, n_13884,
       n_13885;
  wire n_13886, n_13887, n_13888, n_13889, n_13890, n_13891, n_13892,
       n_13893;
  wire n_13894, n_13895, n_13896, n_13897, n_13898, n_13899, n_13900,
       n_13901;
  wire n_13902, n_13903, n_13904, n_13905, n_13906, n_13907, n_13908,
       n_13909;
  wire n_13910, n_13911, n_13912, n_13913, n_13914, n_13915, n_13916,
       n_13917;
  wire n_13918, n_13919, n_13920, n_13921, n_13922, n_13923, n_13924,
       n_13925;
  wire n_13926, n_13927, n_13928, n_13929, n_13930, n_13931, n_13932,
       n_13933;
  wire n_13934, n_13935, n_13936, n_13937, n_13938, n_13939, n_13940,
       n_13942;
  wire n_13943, n_13944, n_13945, n_13946, n_13947, n_13948, n_13949,
       n_13950;
  wire n_13951, n_13952, n_13953, n_13954, n_13955, n_13956, n_13957,
       n_13958;
  wire n_13959, n_13960, n_13961, n_13962, n_13963, n_13964, n_13965,
       n_13966;
  wire n_13967, n_13968, n_13969, n_13970, n_13971, n_13972, n_13973,
       n_13974;
  wire n_13975, n_13976, n_13977, n_13978, n_13979, n_13980, n_13981,
       n_13982;
  wire n_13983, n_13984, n_13985, n_13986, n_13987, n_13988, n_13989,
       n_13990;
  wire n_13991, n_13992, n_13993, n_13994, n_13995, n_13998, n_13999,
       n_14000;
  wire n_14001, n_14002, n_14003, n_14004, n_14005, n_14006, n_14007,
       n_14008;
  wire n_14009, n_14010, n_14011, n_14012, n_14013, n_14014, n_14015,
       n_14016;
  wire n_14017, n_14018, n_14019, n_14020, n_14021, n_14022, n_14023,
       n_14024;
  wire n_14025, n_14026, n_14027, n_14028, n_14029, n_14030, n_14031,
       n_14032;
  wire n_14033, n_14034, n_14035, n_14036, n_14037, n_14038, n_14039,
       n_14040;
  wire n_14041, n_14042, n_14043, n_14044, n_14045, n_14046, n_14047,
       n_14048;
  wire n_14049, n_14050, n_14051, n_14052, n_14053, n_14054, n_14055,
       n_14056;
  wire n_14057, n_14058, n_14059, n_14060, n_14061, n_14062, n_14063,
       n_14064;
  wire n_14065, n_14066, n_14067, n_14068, n_14069, n_14070, n_14071,
       n_14072;
  wire n_14073, n_14074, n_14075, n_14076, n_14077, n_14078, n_14079,
       n_14080;
  wire n_14081, n_14082, n_14083, n_14084, n_14085, n_14086, n_14087,
       n_14088;
  wire n_14089, n_14090, n_14091, n_14092, n_14093, n_14094, n_14095,
       n_14096;
  wire n_14097, n_14098, n_14099, n_14100, n_14101, n_14102, n_14103,
       n_14104;
  wire n_14105, n_14106, n_14107, n_14108, n_14109, n_14110, n_14111,
       n_14112;
  wire n_14113, n_14114, n_14115, n_14116, n_14117, n_14118, n_14119,
       n_14120;
  wire n_14121, n_14122, n_14123, n_14124, n_14125, n_14126, n_14127,
       n_14128;
  wire n_14129, n_14130, n_14131, n_14132, n_14133, n_14134, n_14135,
       n_14136;
  wire n_14137, n_14138, n_14139, n_14140, n_14141, n_14142, n_14143,
       n_14144;
  wire n_14145, n_14146, n_14147, n_14148, n_14149, n_14150, n_14151,
       n_14152;
  wire n_14153, n_14154, n_14155, n_14156, n_14157, n_14158, n_14159,
       n_14160;
  wire n_14161, n_14162, n_14163, n_14164, n_14165, n_14166, n_14167,
       n_14168;
  wire n_14169, n_14170, n_14171, n_14172, n_14173, n_14174, n_14175,
       n_14176;
  wire n_14177, n_14178, n_14179, n_14180, n_14181, n_14182, n_14183,
       n_14184;
  wire n_14185, n_14186, n_14187, n_14188, n_14189, n_14190, n_14191,
       n_14192;
  wire n_14193, n_14194, n_14195, n_14196, n_14197, n_14198, n_14199,
       n_14200;
  wire n_14201, n_14202, n_14203, n_14204, n_14205, n_14206, n_14207,
       n_14208;
  wire n_14209, n_14210, n_14211, n_14212, n_14213, n_14214, n_14215,
       n_14216;
  wire n_14217, n_14218, n_14220, n_14221, n_14222, n_14223, n_14224,
       n_14225;
  wire n_14226, n_14227, n_14228, n_14229, n_14230, n_14231, n_14232,
       n_14233;
  wire n_14234, n_14235, n_14236, n_14237, n_14238, n_14239, n_14240,
       n_14241;
  wire n_14242, n_14243, n_14244, n_14245, n_14246, n_14247, n_14248,
       n_14249;
  wire n_14250, n_14251, n_14252, n_14253, n_14254, n_14255, n_14256,
       n_14257;
  wire n_14258, n_14259, n_14260, n_14261, n_14262, n_14263, n_14264,
       n_14265;
  wire n_14266, n_14267, n_14268, n_14269, n_14270, n_14271, n_14272,
       n_14273;
  wire n_14274, n_14275, n_14276, n_14277, n_14278, n_14279, n_14280,
       n_14281;
  wire n_14282, n_14283, n_14284, n_14285, n_14286, n_14287, n_14288,
       n_14289;
  wire n_14290, n_14291, n_14292, n_14293, n_14294, n_14295, n_14296,
       n_14297;
  wire n_14298, n_14299, n_14300, n_14301, n_14302, n_14303, n_14304,
       n_14305;
  wire n_14306, n_14307, n_14308, n_14309, n_14310, n_14311, n_14312,
       n_14313;
  wire n_14314, n_14315, n_14316, n_14317, n_14318, n_14319, n_14320,
       n_14321;
  wire n_14322, n_14323, n_14324, n_14325, n_14326, n_14327, n_14328,
       n_14329;
  wire n_14330, n_14331, n_14332, n_14333, n_14334, n_14335, n_14336,
       n_14337;
  wire n_14338, n_14339, n_14340, n_14341, n_14342, n_14343, n_14344,
       n_14345;
  wire n_14346, n_14347, n_14348, n_14349, n_14350, n_14351, n_14352,
       n_14353;
  wire n_14354, n_14355, n_14356, n_14357, n_14358, n_14359, n_14360,
       n_14361;
  wire n_14362, n_14363, n_14364, n_14365, n_14366, n_14367, n_14368,
       n_14369;
  wire n_14370, n_14371, n_14372, n_14373, n_14374, n_14375, n_14376,
       n_14377;
  wire n_14378, n_14379, n_14380, n_14381, n_14382, n_14383, n_14384,
       n_14385;
  wire n_14386, n_14387, n_14388, n_14389, n_14390, n_14391, n_14392,
       n_14393;
  wire n_14394, n_14395, n_14396, n_14397, n_14398, n_14399, n_14400,
       n_14401;
  wire n_14402, n_14403, n_14404, n_14405, n_14406, n_14407, n_14408,
       n_14409;
  wire n_14410, n_14411, n_14412, n_14413, n_14414, n_14415, n_14416,
       n_14417;
  wire n_14418, n_14419, n_14420, n_14421, n_14422, n_14423, n_14424,
       n_14425;
  wire n_14426, n_14427, n_14428, n_14429, n_14430, n_14431, n_14432,
       n_14433;
  wire n_14434, n_14435, n_14436, n_14437, n_14438, n_14439, n_14440,
       n_14441;
  wire n_14442, n_14443, n_14444, n_14445, n_14446, n_14447, n_14448,
       n_14449;
  wire n_14450, n_14451, n_14452, n_14453, n_14454, n_14455, n_14456,
       n_14457;
  wire n_14458, n_14459, n_14460, n_14461, n_14462, n_14463, n_14464,
       n_14465;
  wire n_14466, n_14467, n_14468, n_14469, n_14470, n_14471, n_14472,
       n_14473;
  wire n_14474, n_14475, n_14476, n_14477, n_14478, n_14479, n_14480,
       n_14481;
  wire n_14482, n_14483, n_14484, n_14485, n_14486, n_14487, n_14488,
       n_14489;
  wire n_14490, n_14491, n_14492, n_14493, n_14494, n_14495, n_14496,
       n_14497;
  wire n_14498, n_14499, n_14500, n_14501, n_14502, n_14503, n_14504,
       n_14505;
  wire n_14506, n_14507, n_14508, n_14509, n_14510, n_14511, n_14512,
       n_14513;
  wire n_14514, n_14515, n_14516, n_14517, n_14518, n_14519, n_14520,
       n_14521;
  wire n_14522, n_14523, n_14524, n_14525, n_14526, n_14527, n_14528,
       n_14529;
  wire n_14530, n_14531, n_14532, n_14533, n_14534, n_14535, n_14536,
       n_14537;
  wire n_14538, n_14539, n_14540, n_14541, n_14542, n_14543, n_14544,
       n_14545;
  wire n_14546, n_14547, n_14548, n_14549, n_14550, n_14551, n_14552,
       n_14553;
  wire n_14554, n_14555, n_14556, n_14557, n_14558, n_14559, n_14560,
       n_14561;
  wire n_14562, n_14563, n_14564, n_14565, n_14566, n_14567, n_14568,
       n_14569;
  wire n_14570, n_14571, n_14572, n_14573, n_14574, n_14575, n_14576,
       n_14577;
  wire n_14578, n_14582, n_14583, n_14584, n_14585, n_14586, n_14587,
       n_14588;
  wire n_14589, n_14590, n_14591, n_14592, n_14593, n_14594, n_14595,
       n_14596;
  wire n_14597, n_14598, n_14599, n_14600, n_14601, n_14602, n_14603,
       n_14604;
  wire n_14605, n_14606, n_14607, n_14608, n_14609, n_14610, n_14611,
       n_14612;
  wire n_14613, n_14614, n_14615, n_14616, n_14617, n_14618, n_14619,
       n_14620;
  wire n_14621, n_14622, n_14623, n_14624, n_14625, n_14626, n_14627,
       n_14628;
  wire n_14629, n_14630, n_14631, n_14632, n_14633, n_14634, n_14635,
       n_14636;
  wire n_14637, n_14638, n_14639, n_14640, n_14641, n_14642, n_14643,
       n_14644;
  wire n_14645, n_14646, n_14647, n_14648, n_14649, n_14650, n_14651,
       n_14652;
  wire n_14653, n_14654, n_14655, n_14656, n_14657, n_14658, n_14659,
       n_14660;
  wire n_14661, n_14662, n_14663, n_14664, n_14665, n_14666, n_14667,
       n_14668;
  wire n_14669, n_14670, n_14671, n_14672, n_14676, n_14677, n_14678,
       n_14679;
  wire n_14680, n_14681, n_14682, n_14683, n_14684, n_14685, n_14686,
       n_14687;
  wire n_14688, n_14689, n_14690, n_14691, n_14692, n_14693, n_14694,
       n_14695;
  wire n_14696, n_14697, n_14698, n_14699, n_14700, n_14701, n_14702,
       n_14703;
  wire n_14704, n_14705, n_14706, n_14707, n_14708, n_14709, n_14710,
       n_14711;
  wire n_14712, n_14713, n_14714, n_14715, n_14716, n_14717, n_14718,
       n_14719;
  wire n_14720, n_14721, n_14722, n_14723, n_14724, n_14725, n_14726,
       n_14727;
  wire n_14728, n_14729, n_14730, n_14731, n_14732, n_14733, n_14734,
       n_14735;
  wire n_14736, n_14737, n_14738, n_14739, n_14740, n_14741, n_14742,
       n_14743;
  wire n_14744, n_14748, n_14749, n_14750, n_14752, n_14753, n_14754,
       n_14755;
  wire n_14756, n_14757, n_14758, n_14759, n_14760, n_14761, n_14762,
       n_14763;
  wire n_14764, n_14765, n_14766, n_14767, n_14768, n_14769, n_14770,
       n_14771;
  wire n_14772, n_14866, n_14867, n_14871, n_14872, n_14877, n_14879,
       n_14883;
  wire n_14889, n_14896, n_14902, n_14909, n_14910, n_14911, n_14912,
       n_14914;
  wire n_14915, n_14916, n_14917, n_14918, n_14919, n_14920, n_14921,
       n_14922;
  wire n_14924, n_14925, n_14926, n_14927, n_14928, n_14929, n_14930,
       n_14931;
  wire n_14932, n_14933, n_14934, n_14935, n_14937, n_14939, n_14940,
       n_14941;
  wire n_14942, n_14943, n_14944, n_14945, n_14946, n_14947, n_14948,
       n_14950;
  wire n_14951, n_14952, n_14953, n_14954, n_14955, n_14956, n_14957,
       n_14958;
  wire n_14960, n_14961, n_14962, n_14963, n_14964, n_14965, n_14967,
       n_14969;
  wire n_14970, n_14971, n_14972, n_14973, n_14974, n_14975, n_14976,
       n_14977;
  wire n_14978, n_14980, n_14981, n_14982, n_14983, n_14984, n_14985,
       n_14986;
  wire n_14987, n_14989, n_14991, n_14992, n_14993, n_14995, n_14998,
       n_14999;
  wire n_15000, n_15004, n_15005, n_15006, n_15007, n_15008, n_15009,
       n_15010;
  wire n_15012, n_15013, n_15017, n_15019, n_15020, n_15022, n_15023,
       n_15024;
  wire n_15025, n_15026, n_15027, n_15028, n_15029, n_15030, n_15031,
       n_15032;
  wire n_15034, n_15035, n_15037, n_15038, n_15039, n_15041, n_15042,
       n_15043;
  wire n_15045, n_15046, n_15048, n_15050, n_15051, n_15080, n_15090,
       n_15301;
  wire n_15302, n_15304, n_15305, n_15306, n_15308, n_15310, n_15311,
       n_15312;
  wire n_15313, n_15314, n_15315, n_15316, n_15318, n_15319, n_15321,
       n_15323;
  wire n_15324, n_15326, n_15328, n_15329, n_15330, n_15331, n_15333,
       n_15334;
  wire n_15335, n_15336, n_15337, n_15338, n_15339, n_15340, n_15342,
       n_15344;
  wire n_15345, n_15346, n_15347, n_15349, n_15351, n_15353, n_15355,
       n_15357;
  wire n_15359, n_15361, n_15362, n_15363, n_15364, n_15366, n_15368,
       n_15370;
  wire n_15372, n_15373, n_15374, n_15375, n_15376, n_15377, n_15379,
       n_15381;
  wire n_15383, n_15385, n_15386, n_15387, n_15388, n_15389, n_15391,
       n_15392;
  wire n_15394, n_15396, n_15397, n_15398, n_15400, n_15401, n_15404,
       n_15405;
  wire n_15408, n_15409, n_15410, n_15411, n_15413, n_15414, n_15415,
       n_15417;
  wire n_15418, n_15420, n_15421, n_15423, n_15424, n_15427, n_15429,
       n_15430;
  wire n_15431, n_15432, n_15433, n_15434, n_15435, n_15436, n_15439,
       n_15440;
  wire n_15442, n_15443, n_15444, n_15445, n_15446, n_15447, n_15448,
       n_15449;
  wire n_15450, n_15451, n_15452, n_15453, n_15454, n_15455, n_15456,
       n_15457;
  wire n_15458, n_15459, n_15460, n_15461, n_15462, n_15463, n_15464,
       n_15465;
  wire n_15466, n_15467, n_15468, n_15469, n_15470, n_15471, n_15472,
       n_15473;
  wire n_15474, n_15475, n_15476, n_15477, n_15478, n_15479, n_15480,
       n_15481;
  wire n_15482, n_15483, n_15484, n_15485, n_15486, n_15487, n_15488,
       n_15489;
  wire n_15490, n_15491, n_15492, n_15493, n_15494, n_15495, n_15496,
       n_15497;
  wire n_15498, n_15499, n_15500, n_15501, n_15502, n_15503, n_15504,
       n_15505;
  wire n_15506, n_15507, n_15508, n_15509, n_15510, n_15511, n_15512,
       n_15513;
  wire n_15514, n_15515, n_15516, n_15517, n_15518, n_15519, n_15526,
       n_15527;
  wire n_15528, n_15531, n_15538, n_15539, n_15540, n_15545, n_15546,
       n_15549;
  wire n_15552, n_15573, n_15574, n_15575, n_15576, n_15577, n_15578,
       n_15579;
  wire n_15580, n_15581, n_15582, n_15585, n_15588, n_15591, n_15594,
       n_15597;
  wire n_15600, n_15605, n_15606, n_15611, n_15612, n_15615, n_15618,
       n_15621;
  wire n_15624, n_15627, n_15630, n_15633, n_15636, n_15639, n_15646,
       n_15647;
  wire n_15648, n_15651, n_15656, n_15657, n_15660, n_15663, n_15666,
       n_15669;
  wire n_15672, n_15675, n_15678, n_15681, n_15686, n_15687, n_15690,
       n_15695;
  wire n_15696, n_15703, n_15704, n_15705, n_15708, n_15711, n_15714,
       n_15717;
  wire n_15724, n_15725, n_15726, n_15729, n_15738, n_15739, n_15740,
       n_15741;
  wire n_15750, n_15751, n_15752, n_15753, n_15762, n_15763, n_15764,
       n_15765;
  wire n_15774, n_15775, n_15776, n_15777, n_15786, n_15787, n_15788,
       n_15789;
  wire n_15798, n_15799, n_15800, n_15801, n_15804, n_15819, n_15820,
       n_15821;
  wire n_15822, n_15823, n_15824, n_15825, n_15840, n_15841, n_15842,
       n_15843;
  wire n_15844, n_15845, n_15846, n_15861, n_15862, n_15863, n_15864,
       n_15865;
  wire n_15866, n_15867, n_15882, n_15883, n_15884, n_15885, n_15886,
       n_15887;
  wire n_15888, n_15903, n_15904, n_15905, n_15906, n_15907, n_15908,
       n_15909;
  wire n_15924, n_15925, n_15926, n_15927, n_15928, n_15929, n_15930,
       n_15943;
  wire n_15944, n_15945, n_15946, n_15947, n_15948, n_15951, n_15954,
       n_15957;
  wire n_15960, n_15963, n_15966, n_15975, n_15976, n_15977, n_15978,
       n_15985;
  wire n_15986, n_15987, n_15990, n_15997, n_15998, n_15999, n_16006,
       n_16007;
  wire n_16008, n_16023, n_16024, n_16025, n_16026, n_16027, n_16028,
       n_16029;
  wire n_16032, n_16043, n_16044, n_16045, n_16046, n_16047, n_16056,
       n_16057;
  wire n_16058, n_16059, n_16068, n_16069, n_16070, n_16071, n_16080,
       n_16081;
  wire n_16082, n_16083, n_16086, n_16089, n_16092, n_16099, n_16100,
       n_16101;
  wire n_16106, n_16107, n_16110, n_16124, n_16125, n_16139, n_16140,
       n_16143;
  wire n_16148, n_16149, n_16152, n_16155, n_16158, n_16165, n_16166,
       n_16167;
  wire n_16170, n_16182, n_16183, n_16184, n_16185, n_16190, n_16191,
       n_16196;
  wire n_16197, n_16206, n_16207, n_16208, n_16209, n_16214, n_16215,
       n_16220;
  wire n_16221, n_16224, n_16227, n_16232, n_16233, n_16247, n_16248,
       n_16262;
  wire n_16263, n_16270, n_16271, n_16272, n_16279, n_16280, n_16284,
       n_16287;
  wire n_16290, n_16299, n_16300, n_16301, n_16302, n_16311, n_16312,
       n_16313;
  wire n_16314, n_16317, n_16322, n_16323, n_16328, n_16329, n_16332,
       n_16337;
  wire n_16343, n_16344, n_16349, n_16350, n_16353, n_16356, n_16361,
       n_16362;
  wire n_16367, n_16368, n_16373, n_16374, n_16379, n_16380, n_16385,
       n_16386;
  wire n_16395, n_16396, n_16397, n_16398, n_16407, n_16408, n_16409,
       n_16410;
  wire n_16415, n_16416, n_16421, n_16422, n_16427, n_16428, n_16433,
       n_16434;
  wire n_16439, n_16440, n_16443, n_16446, n_16451, n_16452, n_16455,
       n_16458;
  wire n_16461, n_16464, n_16467, n_16472, n_16473, n_16478, n_16479,
       n_16484;
  wire n_16485, n_16490, n_16491, n_16496, n_16497, n_16502, n_16503,
       n_16508;
  wire n_16509, n_16514, n_16515, n_16520, n_16521, n_16526, n_16527,
       n_16532;
  wire n_16533, n_16538, n_16539, n_16544, n_16545, n_16550, n_16551,
       n_16556;
  wire n_16557, n_16562, n_16563, n_16568, n_16569, n_16574, n_16575,
       n_16580;
  wire n_16581, n_16586, n_16587, n_16592, n_16593, n_16598, n_16599,
       n_16604;
  wire n_16605, n_16610, n_16611, n_16616, n_16617, n_16622, n_16623,
       n_16628;
  wire n_16629, n_16634, n_16635, n_16640, n_16641, n_16646, n_16647,
       n_16652;
  wire n_16653, n_16658, n_16659, n_16664, n_16665, n_16670, n_16671,
       n_16676;
  wire n_16677, n_16682, n_16683, n_16688, n_16689, n_16694, n_16695,
       n_16700;
  wire n_16701, n_16706, n_16707, n_16712, n_16713, n_16718, n_16719,
       n_16724;
  wire n_16725, n_16730, n_16731, n_16736, n_16737, n_16742, n_16743,
       n_16748;
  wire n_16749, n_16754, n_16755, n_16760, n_16761, n_16766, n_16767,
       n_16772;
  wire n_16773, n_16778, n_16779, n_16784, n_16785, n_16790, n_16791,
       n_16796;
  wire n_16797, n_16802, n_16803, n_16808, n_16809, n_16814, n_16815,
       n_16820;
  wire n_16821, n_16826, n_16827, n_16832, n_16833, n_16838, n_16839,
       n_16844;
  wire n_16845, n_16850, n_16851, n_16856, n_16857, n_16862, n_16863,
       n_16868;
  wire n_16869, n_16874, n_16875, n_16880, n_16881, n_16886, n_16887,
       n_16892;
  wire n_16893, n_16898, n_16899, n_16904, n_16905, n_16910, n_16911,
       n_16916;
  wire n_16917, n_16922, n_16923, n_16928, n_16929, n_16934, n_16935,
       n_16940;
  wire n_16941, n_16946, n_16947, n_16952, n_16953, n_16958, n_16959,
       n_16964;
  wire n_16965, n_16970, n_16971, n_16976, n_16977, n_16982, n_16983,
       n_16988;
  wire n_16989, n_16994, n_16995, n_17000, n_17001, n_17006, n_17007,
       n_17012;
  wire n_17013, n_17018, n_17019, n_17024, n_17025, n_17030, n_17031,
       n_17036;
  wire n_17037, n_17042, n_17043, n_17072, n_17073, n_17074, n_17075,
       n_17076;
  wire n_17077, n_17078, n_17079, n_17080, n_17081, n_17082, n_17083,
       n_17084;
  wire n_17085, n_17118, n_17119, n_17120, n_17121, n_17122, n_17123,
       n_17124;
  wire n_17125, n_17126, n_17127, n_17128, n_17129, n_17130, n_17131,
       n_17132;
  wire n_17133, n_17166, n_17167, n_17168, n_17169, n_17170, n_17171,
       n_17172;
  wire n_17173, n_17174, n_17175, n_17176, n_17177, n_17178, n_17179,
       n_17180;
  wire n_17181, n_17214, n_17215, n_17216, n_17217, n_17218, n_17219,
       n_17220;
  wire n_17221, n_17222, n_17223, n_17224, n_17225, n_17226, n_17227,
       n_17228;
  wire n_17229, n_17262, n_17263, n_17264, n_17265, n_17266, n_17267,
       n_17268;
  wire n_17269, n_17270, n_17271, n_17272, n_17273, n_17274, n_17275,
       n_17276;
  wire n_17277, n_17310, n_17311, n_17312, n_17313, n_17314, n_17315,
       n_17316;
  wire n_17317, n_17318, n_17319, n_17320, n_17321, n_17322, n_17323,
       n_17324;
  wire n_17325, n_17358, n_17359, n_17360, n_17361, n_17362, n_17363,
       n_17364;
  wire n_17365, n_17366, n_17367, n_17368, n_17369, n_17370, n_17371,
       n_17372;
  wire n_17373, n_17406, n_17407, n_17408, n_17409, n_17410, n_17411,
       n_17412;
  wire n_17413, n_17414, n_17415, n_17416, n_17417, n_17418, n_17419,
       n_17420;
  wire n_17421, n_17454, n_17455, n_17456, n_17457, n_17458, n_17459,
       n_17460;
  wire n_17461, n_17462, n_17463, n_17464, n_17465, n_17466, n_17467,
       n_17468;
  wire n_17469, n_17502, n_17503, n_17504, n_17505, n_17506, n_17507,
       n_17508;
  wire n_17509, n_17510, n_17511, n_17512, n_17513, n_17514, n_17515,
       n_17516;
  wire n_17517, n_17550, n_17551, n_17552, n_17553, n_17554, n_17555,
       n_17556;
  wire n_17557, n_17558, n_17559, n_17560, n_17561, n_17562, n_17563,
       n_17564;
  wire n_17565, n_17598, n_17599, n_17600, n_17601, n_17602, n_17603,
       n_17604;
  wire n_17605, n_17606, n_17607, n_17608, n_17609, n_17610, n_17611,
       n_17612;
  wire n_17613, n_17646, n_17647, n_17648, n_17649, n_17650, n_17651,
       n_17652;
  wire n_17653, n_17654, n_17655, n_17656, n_17657, n_17658, n_17659,
       n_17660;
  wire n_17661, n_17694, n_17695, n_17696, n_17697, n_17698, n_17699,
       n_17700;
  wire n_17701, n_17702, n_17703, n_17704, n_17705, n_17706, n_17707,
       n_17708;
  wire n_17709, n_17742, n_17743, n_17744, n_17745, n_17746, n_17747,
       n_17748;
  wire n_17749, n_17750, n_17751, n_17752, n_17753, n_17754, n_17755,
       n_17756;
  wire n_17757, n_17790, n_17791, n_17792, n_17793, n_17794, n_17795,
       n_17796;
  wire n_17797, n_17798, n_17799, n_17800, n_17801, n_17802, n_17803,
       n_17804;
  wire n_17805, n_17838, n_17839, n_17840, n_17841, n_17842, n_17843,
       n_17844;
  wire n_17845, n_17846, n_17847, n_17848, n_17849, n_17850, n_17851,
       n_17852;
  wire n_17853, n_17886, n_17887, n_17888, n_17889, n_17890, n_17891,
       n_17892;
  wire n_17893, n_17894, n_17895, n_17896, n_17897, n_17898, n_17899,
       n_17900;
  wire n_17901, n_17934, n_17935, n_17936, n_17937, n_17938, n_17939,
       n_17940;
  wire n_17941, n_17942, n_17943, n_17944, n_17945, n_17946, n_17947,
       n_17948;
  wire n_17949, n_17982, n_17983, n_17984, n_17985, n_17986, n_17987,
       n_17988;
  wire n_17989, n_17990, n_17991, n_17992, n_17993, n_17994, n_17995,
       n_17996;
  wire n_17997, n_18030, n_18031, n_18032, n_18033, n_18034, n_18035,
       n_18036;
  wire n_18037, n_18038, n_18039, n_18040, n_18041, n_18042, n_18043,
       n_18044;
  wire n_18045, n_18078, n_18079, n_18080, n_18081, n_18082, n_18083,
       n_18084;
  wire n_18085, n_18086, n_18087, n_18088, n_18089, n_18090, n_18091,
       n_18092;
  wire n_18093, n_18098, n_18104, n_18110, n_18116, n_18122, n_18123,
       n_18140;
  wire n_18141, n_18146, n_18147, n_18152, n_18153, n_18158, n_18159,
       n_18164;
  wire n_18165, n_18170, n_18171, n_18176, n_18177, n_18182, n_18183,
       n_18188;
  wire n_18189, n_18194, n_18195, n_18200, n_18201, n_18206, n_18214,
       n_18215;
  wire n_18216, n_18221, n_18233, n_18234, n_18235, n_18236, n_18237,
       n_18242;
  wire n_18243, n_18254, n_18255, n_18256, n_18257, n_18258, n_18269,
       n_18270;
  wire n_18271, n_18272, n_18273, n_18284, n_18285, n_18286, n_18287,
       n_18288;
  wire n_18299, n_18300, n_18301, n_18302, n_18303, n_18308, n_18309,
       n_18314;
  wire n_18315, n_18322, n_18324, n_18331, n_18332, n_18333, n_18338,
       n_18339;
  wire n_18344, n_18345, n_18350, n_18351, n_18358, n_18359, n_18360,
       n_18371;
  wire n_18372, n_18373, n_18374, n_18375, n_18386, n_18387, n_18388,
       n_18389;
  wire n_18390, n_18401, n_18402, n_18403, n_18404, n_18405, n_18410,
       n_18411;
  wire n_18416, n_18417, n_18422, n_18423, n_18428, n_18429, n_18434,
       n_18435;
  wire n_18440, n_18441, n_18446, n_18452, n_18458, n_18470, n_18471,
       n_18472;
  wire n_18473, n_18474, n_18485, n_18486, n_18487, n_18488, n_18489,
       n_18494;
  wire n_18495, n_18500, n_18501, n_18506, n_18507, n_18512, n_18518,
       n_18519;
  wire n_18526, n_18527, n_18528, n_18535, n_18536, n_18537, n_18542,
       n_18543;
  wire n_18548, n_18549, n_18554, n_18555, n_18560, n_18561, n_18566,
       n_18567;
  wire n_18572, n_18573, n_18578, n_18579, n_18584, n_18585, n_18590,
       n_18591;
  wire n_18596, n_18597, n_18602, n_18610, n_18611, n_18612, n_18617,
       n_18623;
  wire n_18624, n_18629, n_18635, n_18641, n_18653, n_18654, n_18655,
       n_18656;
  wire n_18657, n_18668, n_18669, n_18670, n_18671, n_18672, n_18677,
       n_18678;
  wire n_18683, n_18684, n_18691, n_18693, n_18698, n_18699, n_18713,
       n_18714;
  wire n_18719, n_18720, n_18725, n_18731, n_18732, n_18737, n_18738,
       n_18743;
  wire n_18744, n_18747, n_18750, n_18755, n_18756, n_18761, n_18762,
       n_18767;
  wire n_18768, n_18773, n_18774, n_18779, n_18780, n_18785, n_18786,
       n_18797;
  wire n_18798, n_18799, n_18800, n_18801, n_18806, n_18807, n_18812,
       n_18813;
  wire n_18818, n_18819, n_18824, n_18825, n_18830, n_18836, n_18842,
       n_18843;
  wire n_18848, n_18849, n_18854, n_18858, n_18861, n_18866, n_18867,
       n_18872;
  wire n_18873, n_18878, n_18879, n_18895, n_18896, n_18897, n_18902,
       n_18903;
  wire n_18908, n_18914, n_18920, n_18921, n_18926, n_18927, n_18932,
       n_18933;
  wire n_18938, n_18939, n_18944, n_18945, n_18950, n_18951, n_18956,
       n_18957;
  wire n_18962, n_18963, n_18968, n_18969, n_18974, n_18975, n_18980,
       n_18981;
  wire n_18986, n_18987, n_18992, n_18993, n_18998, n_19004, n_19005,
       n_19010;
  wire n_19011, n_19016, n_19026, n_19027, n_19028, n_19029, n_19032,
       n_19035;
  wire n_19048, n_19050, n_19051, n_19052, n_19053, n_19058, n_19059,
       n_19064;
  wire n_19065, n_19070, n_19071, n_19074, n_19079, n_19080, n_19087,
       n_19088;
  wire n_19089, n_19103, n_19104, n_19109, n_19110, n_19115, n_19116,
       n_19123;
  wire n_19124, n_19125, n_19130, n_19131, n_19138, n_19139, n_19140,
       n_19153;
  wire n_19154, n_19155, n_19156, n_19157, n_19158, n_19161, n_19166,
       n_19167;
  wire n_19170, n_19175, n_19176, n_19181, n_19182, n_19187, n_19193,
       n_19199;
  wire n_19205, n_19211, n_19212, n_19217, n_19218, n_19223, n_19224,
       n_19233;
  wire n_19234, n_19235, n_19236, n_19241, n_19242, n_19247, n_19248,
       n_19253;
  wire n_19254, n_19259, n_19260, n_19265, n_19266, n_19271, n_19272,
       n_19277;
  wire n_19278, n_19283, n_19284, n_19289, n_19290, n_19293, n_19296,
       n_19299;
  wire n_19304, n_19305, n_19308, n_19313, n_19314, n_19319, n_19320,
       n_19325;
  wire n_19326, n_19337, n_19338, n_19339, n_19340, n_19341, n_19346,
       n_19347;
  wire n_19352, n_19353, n_19364, n_19365, n_19366, n_19367, n_19368,
       n_19373;
  wire n_19374, n_19379, n_19380, n_19391, n_19392, n_19393, n_19394,
       n_19395;
  wire n_19416, n_19417, n_19418, n_19419, n_19420, n_19421, n_19422,
       n_19423;
  wire n_19424, n_19425, n_19430, n_19431, n_19436, n_19437, n_19442,
       n_19443;
  wire n_19448, n_19449, n_19454, n_19455, n_19460, n_19461, n_19466,
       n_19467;
  wire n_19472, n_19473, n_19478, n_19479, n_19484, n_19485, n_19492,
       n_19493;
  wire n_19494, n_19502, n_19510, n_19511, n_19512, n_19515, n_19518,
       n_19523;
  wire n_19524, n_19527, n_19532, n_19533, n_19538, n_19539, n_19544,
       n_19545;
  wire n_19562, n_19563, n_19564, n_19565, n_19566, n_19567, n_19568,
       n_19569;
  wire n_19572, n_19575, n_19580, n_19581, n_19586, n_19587, n_19592,
       n_19593;
  wire n_19600, n_19601, n_19602, n_19607, n_19608, n_19615, n_19616,
       n_19617;
  wire n_19620, n_19623, n_19626, n_19635, n_19636, n_19637, n_19638,
       n_19643;
  wire n_19644, n_19649, n_19650, n_19655, n_19656, n_19661, n_19662,
       n_19667;
  wire n_19668, n_19673, n_19674, n_19679, n_19680, n_19685, n_19686,
       n_19691;
  wire n_19692, n_19697, n_19698, n_19715, n_19716, n_19717, n_19718,
       n_19719;
  wire n_19720, n_19721, n_19722, n_19725, n_19730, n_19731, n_19742,
       n_19743;
  wire n_19744, n_19745, n_19746, n_19749, n_19760, n_19761, n_19762,
       n_19763;
  wire n_19764, n_19769, n_19770, n_19775, n_19776, n_19779, n_19786,
       n_19787;
  wire n_19788, n_19795, n_19796, n_19797, n_19800, n_19803, n_19808,
       n_19809;
  wire n_19818, n_19819, n_19820, n_19821, n_19826, n_19827, n_19832,
       n_19833;
  wire n_19838, n_19839, n_19844, n_19845, n_19850, n_19851, n_19856,
       n_19857;
  wire n_19862, n_19863, n_19868, n_19869, n_19872, n_19875, n_19880,
       n_19881;
  wire n_19886, n_19887, n_19898, n_19899, n_19900, n_19901, n_19902,
       n_19907;
  wire n_19908, n_19915, n_19917, n_19922, n_19923, n_19940, n_19941,
       n_19942;
  wire n_19943, n_19944, n_19945, n_19946, n_19947, n_19950, n_19953,
       n_19964;
  wire n_19965, n_19966, n_19967, n_19968, n_19973, n_19974, n_19977,
       n_19982;
  wire n_19983, n_19986, n_19989, n_19992, n_20001, n_20002, n_20003,
       n_20004;
  wire n_20009, n_20010, n_20015, n_20016, n_20021, n_20022, n_20027,
       n_20028;
  wire n_20033, n_20034, n_20039, n_20040, n_20045, n_20046, n_20051,
       n_20052;
  wire n_20059, n_20061, n_20064, n_20067, n_20072, n_20073, n_20094,
       n_20095;
  wire n_20096, n_20097, n_20098, n_20099, n_20100, n_20101, n_20102,
       n_20103;
  wire n_20108, n_20109, n_20114, n_20115, n_20120, n_20121, n_20126,
       n_20127;
  wire n_20132, n_20133, n_20138, n_20139, n_20144, n_20145, n_20150,
       n_20151;
  wire n_20168, n_20169, n_20170, n_20171, n_20172, n_20173, n_20174,
       n_20175;
  wire n_20178, n_20183, n_20184, n_20187, n_20190, n_20199, n_20200,
       n_20201;
  wire n_20202, n_20207, n_20208, n_20213, n_20214, n_20219, n_20220,
       n_20225;
  wire n_20226, n_20231, n_20232, n_20237, n_20238, n_20243, n_20244,
       n_20249;
  wire n_20250, n_20255, n_20256, n_20259, n_20268, n_20269, n_20270,
       n_20271;
  wire n_20288, n_20289, n_20290, n_20291, n_20292, n_20293, n_20294,
       n_20295;
  wire n_20300, n_20301, n_20304, n_20309, n_20310, n_20313, n_20324,
       n_20325;
  wire n_20326, n_20327, n_20328, n_20335, n_20336, n_20337, n_20342,
       n_20343;
  wire n_20348, n_20349, n_20354, n_20355, n_20360, n_20361, n_20366,
       n_20367;
  wire n_20372, n_20373, n_20378, n_20379, n_20384, n_20385, n_20390,
       n_20391;
  wire n_20396, n_20397, n_20402, n_20403, n_20408, n_20409, n_20414,
       n_20415;
  wire n_20420, n_20421, n_20426, n_20427, n_20432, n_20433, n_20436,
       n_20439;
  wire n_20442, n_20445, n_20448, n_20451, n_20454, n_20457, n_20460,
       n_20463;
  wire n_20466, n_20469, n_20472, n_20475, n_20478, n_20481, n_20484,
       n_20487;
  wire n_20490, n_20493, n_20496, n_20499, n_20502, n_20505, n_20508,
       n_20511;
  wire n_20514, n_20517, n_20520, n_20523, n_20526, n_20529, n_20532,
       n_20539;
  wire n_20540, n_20541, n_20548, n_20549, n_20550, n_20555, n_20556,
       n_20561;
  wire n_20562, n_20567, n_20568, n_20573, n_20574, n_20579, n_20580,
       n_20585;
  wire n_20586, n_20591, n_20592, n_20597, n_20598, n_20603, n_20604,
       n_20609;
  wire n_20610, n_20615, n_20616, n_20621, n_20622, n_20627, n_20628,
       n_20633;
  wire n_20634, n_20639, n_20640, n_20645, n_20646, n_20653, n_20654,
       n_20655;
  wire n_20660, n_20661, n_20666, n_20667, n_20672, n_20673, n_20678,
       n_20679;
  wire n_20684, n_20685, n_20690, n_20691, n_20696, n_20697, n_20702,
       n_20703;
  wire n_20708, n_20709, n_20714, n_20715, n_20720, n_20721, n_20726,
       n_20727;
  wire n_20732, n_20733, n_20738, n_20739, n_20744, n_20745, n_20750,
       n_20751;
  wire n_20756, n_20757, n_20762, n_20763, n_20768, n_20769, n_20774,
       n_20775;
  wire n_20780, n_20781, n_20786, n_20787, n_20792, n_20793, n_20798,
       n_20799;
  wire n_20802, n_20805, n_20808, n_20811, n_20814, n_20817, n_20820,
       n_20823;
  wire n_20826, n_20829, n_20832, n_20835, n_20838, n_20841, n_20844,
       n_20847;
  wire n_20850, n_20853, n_20856, n_20859, n_20862, n_20865, n_20868,
       n_20871;
  wire n_20874, n_20877, n_20880, n_20883, n_20886, n_20889, n_20892,
       n_20895;
  wire n_20898, n_20901, n_20904, n_20907, n_20910, n_20913, n_20916,
       n_20919;
  wire n_20922, n_20925, n_20928, n_20931, n_20934, n_20937, n_20940,
       n_20943;
  wire n_20946, n_20949, n_20952, n_20955, n_20958, n_20961, n_20964,
       n_20967;
  wire n_20970, n_20973, n_20976, n_20979, n_20982, n_20985, n_20988,
       n_20991;
  wire n_20994, n_20997, n_21000, n_21003, n_21006, n_21009, n_21012,
       n_21015;
  wire n_21018, n_21023, n_21024, n_21029, n_21030, n_21843, n_21844,
       n_21845;
  wire n_21846, n_21847, n_21848, n_21849, n_21850, n_21851, n_21852,
       n_21853;
  wire n_21854, n_21855, n_21856, n_21857, n_21858, n_21859, n_21860,
       n_21861;
  wire n_21862, n_21863, n_21864, n_21865, n_21866, n_21867, n_21868,
       n_21869;
  wire n_21870, n_21871, n_21872, n_21873, n_21874, n_21877, n_21878,
       n_21879;
  wire n_21880, n_21881, n_21882, n_21883, n_21884, n_21885, n_21886,
       n_21887;
  wire n_21888, n_21891, n_21892, n_21893, n_21894, n_21895, n_21896,
       n_21897;
  wire n_21898, n_21899, n_21900, n_21901, n_21902, n_21905, n_21906,
       n_21907;
  wire n_21908, n_21909, n_21910, n_21911, n_21912, n_21913, n_21914,
       n_21915;
  wire n_21916, n_21917, n_21918, n_21919, n_21920, n_21921, n_21922,
       n_21923;
  wire n_21924, n_21925, n_21926, n_21927, n_21928, n_21929, n_21930,
       n_21931;
  wire n_21932, n_21933, n_21934, n_21935, n_21936, n_21937, n_21938,
       n_21939;
  wire n_21940, n_21941, n_21942, n_21945, n_21946, n_21947, n_21948,
       n_21949;
  wire n_21950, n_21951, n_21952, n_21953, n_21954, n_21955, n_21956,
       n_21957;
  wire n_21958, n_21959, n_21960, n_21961, n_21962, n_21963, n_21964,
       n_21965;
  wire n_21966, n_21967, n_21968, n_21969, n_21970, n_21971, n_21972,
       n_21973;
  wire n_21974, n_21975, n_21976, n_21977, n_21978, n_21979, n_21980,
       n_21981;
  wire n_21982, n_21983, n_21984, n_21985, n_21986, n_21987, n_21988,
       n_21989;
  wire n_21990, n_21991, n_21992, n_21993, n_21994, n_21995, n_21996,
       n_21997;
  wire n_21998, n_21999, n_22000, n_22001, n_22002, n_22003, n_22004,
       n_22005;
  wire n_22006, n_22007, n_22008, n_22009, n_22010, n_22011, n_22012,
       n_22013;
  wire n_22014, n_22015, n_22016, n_22017, n_22018, n_22019, n_22020,
       n_22021;
  wire n_22022, n_22023, n_22024, n_22025, n_22026, n_22027, n_22028,
       n_22029;
  wire n_22030, n_22031, n_22032, n_22033, n_22034, n_22035, n_22036,
       n_22037;
  wire n_22038, n_22039, n_22040, n_22041, n_22042, n_22043, n_22044,
       n_22045;
  wire n_22046, n_22047, n_22048, n_22049, n_22050, n_22051, n_22052,
       n_22053;
  wire n_22054, n_22055, n_22056, n_22057, n_22058, n_22059, n_22060,
       n_22061;
  wire n_22062, n_22063, n_22064, n_22065, n_22066, n_22067, n_22068,
       n_22069;
  wire n_22070, n_22071, n_22072, n_22073, n_22074, n_22075, n_22077,
       n_22078;
  wire n_22079, n_22080, n_22081, n_22082, n_22083, n_22084, n_22085,
       n_22086;
  wire n_22087, n_22088, n_22089, n_22090, n_22091, n_22092, n_22093,
       n_22094;
  wire n_22095, n_22096, n_22097, n_22098, n_22099;
  CDN_flop \data_stack_mem_reg[0][0] (.clk (clk), .d (n_14646), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [0]));
  CDN_flop \data_stack_mem_reg[0][1] (.clk (clk), .d (n_14647), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [1]));
  CDN_flop \data_stack_mem_reg[0][2] (.clk (clk), .d (n_14648), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [2]));
  CDN_flop \data_stack_mem_reg[0][3] (.clk (clk), .d (n_14649), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [3]));
  CDN_flop \data_stack_mem_reg[0][4] (.clk (clk), .d (n_14643), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [4]));
  CDN_flop \data_stack_mem_reg[0][5] (.clk (clk), .d (n_14645), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [5]));
  CDN_flop \data_stack_mem_reg[0][6] (.clk (clk), .d (n_14642), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [6]));
  CDN_flop \data_stack_mem_reg[0][7] (.clk (clk), .d (n_14644), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [7]));
  CDN_flop \data_stack_mem_reg[1][0] (.clk (clk), .d (n_14639), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [0]));
  CDN_flop \data_stack_mem_reg[1][1] (.clk (clk), .d (n_14638), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [1]));
  CDN_flop \data_stack_mem_reg[1][2] (.clk (clk), .d (n_14637), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [2]));
  CDN_flop \data_stack_mem_reg[1][3] (.clk (clk), .d (n_14636), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [3]));
  CDN_flop \data_stack_mem_reg[1][4] (.clk (clk), .d (n_14635), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [4]));
  CDN_flop \data_stack_mem_reg[1][5] (.clk (clk), .d (n_14634), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [5]));
  CDN_flop \data_stack_mem_reg[1][6] (.clk (clk), .d (n_14633), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [6]));
  CDN_flop \data_stack_mem_reg[1][7] (.clk (clk), .d (n_14632), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [7]));
  CDN_flop \data_stack_mem_reg[2][0] (.clk (clk), .d (n_14595), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [0]));
  CDN_flop \data_stack_mem_reg[2][1] (.clk (clk), .d (n_14594), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [1]));
  CDN_flop \data_stack_mem_reg[2][2] (.clk (clk), .d (n_14593), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [2]));
  CDN_flop \data_stack_mem_reg[2][3] (.clk (clk), .d (n_14592), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [3]));
  CDN_flop \data_stack_mem_reg[2][4] (.clk (clk), .d (n_14589), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [4]));
  CDN_flop \data_stack_mem_reg[2][5] (.clk (clk), .d (n_14590), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [5]));
  CDN_flop \data_stack_mem_reg[2][6] (.clk (clk), .d (n_14591), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [6]));
  CDN_flop \data_stack_mem_reg[2][7] (.clk (clk), .d (n_14596), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [7]));
  CDN_flop \data_stack_mem_reg[3][0] (.clk (clk), .d (n_14600), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [0]));
  CDN_flop \data_stack_mem_reg[3][1] (.clk (clk), .d (n_14604), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [1]));
  CDN_flop \data_stack_mem_reg[3][2] (.clk (clk), .d (n_14605), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [2]));
  CDN_flop \data_stack_mem_reg[3][3] (.clk (clk), .d (n_14601), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [3]));
  CDN_flop \data_stack_mem_reg[3][4] (.clk (clk), .d (n_14602), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [4]));
  CDN_flop \data_stack_mem_reg[3][5] (.clk (clk), .d (n_14606), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [5]));
  CDN_flop \data_stack_mem_reg[3][6] (.clk (clk), .d (n_14599), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [6]));
  CDN_flop \data_stack_mem_reg[3][7] (.clk (clk), .d (n_14603), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [7]));
  CDN_flop \data_stack_mem_reg[4][0] (.clk (clk), .d (n_14654), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [0]));
  CDN_flop \data_stack_mem_reg[4][1] (.clk (clk), .d (n_14660), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [1]));
  CDN_flop \data_stack_mem_reg[4][2] (.clk (clk), .d (n_14653), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [2]));
  CDN_flop \data_stack_mem_reg[4][3] (.clk (clk), .d (n_14659), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [3]));
  CDN_flop \data_stack_mem_reg[4][4] (.clk (clk), .d (n_14658), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [4]));
  CDN_flop \data_stack_mem_reg[4][5] (.clk (clk), .d (n_14657), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [5]));
  CDN_flop \data_stack_mem_reg[4][6] (.clk (clk), .d (n_14656), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [6]));
  CDN_flop \data_stack_mem_reg[4][7] (.clk (clk), .d (n_14655), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [7]));
  CDN_flop \data_stack_mem_reg[5][0] (.clk (clk), .d (n_14692), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [0]));
  CDN_flop \data_stack_mem_reg[5][1] (.clk (clk), .d (n_14690), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [1]));
  CDN_flop \data_stack_mem_reg[5][2] (.clk (clk), .d (n_14691), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [2]));
  CDN_flop \data_stack_mem_reg[5][3] (.clk (clk), .d (n_14689), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [3]));
  CDN_flop \data_stack_mem_reg[5][4] (.clk (clk), .d (n_14688), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [4]));
  CDN_flop \data_stack_mem_reg[5][5] (.clk (clk), .d (n_14687), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [5]));
  CDN_flop \data_stack_mem_reg[5][6] (.clk (clk), .d (n_14686), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [6]));
  CDN_flop \data_stack_mem_reg[5][7] (.clk (clk), .d (n_14685), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [7]));
  CDN_flop \data_stack_mem_reg[6][0] (.clk (clk), .d (n_14621), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [0]));
  CDN_flop \data_stack_mem_reg[6][1] (.clk (clk), .d (n_14622), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [1]));
  CDN_flop \data_stack_mem_reg[6][2] (.clk (clk), .d (n_14623), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [2]));
  CDN_flop \data_stack_mem_reg[6][3] (.clk (clk), .d (n_14624), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [3]));
  CDN_flop \data_stack_mem_reg[6][4] (.clk (clk), .d (n_14625), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [4]));
  CDN_flop \data_stack_mem_reg[6][5] (.clk (clk), .d (n_14626), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [5]));
  CDN_flop \data_stack_mem_reg[6][6] (.clk (clk), .d (n_14627), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [6]));
  CDN_flop \data_stack_mem_reg[6][7] (.clk (clk), .d (n_14628), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [7]));
  CDN_flop \data_stack_mem_reg[7][0] (.clk (clk), .d (n_14612), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [0]));
  CDN_flop \data_stack_mem_reg[7][1] (.clk (clk), .d (n_14614), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [1]));
  CDN_flop \data_stack_mem_reg[7][2] (.clk (clk), .d (n_14615), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [2]));
  CDN_flop \data_stack_mem_reg[7][3] (.clk (clk), .d (n_14617), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [3]));
  CDN_flop \data_stack_mem_reg[7][4] (.clk (clk), .d (n_14616), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [4]));
  CDN_flop \data_stack_mem_reg[7][5] (.clk (clk), .d (n_14611), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [5]));
  CDN_flop \data_stack_mem_reg[7][6] (.clk (clk), .d (n_14618), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [6]));
  CDN_flop \data_stack_mem_reg[7][7] (.clk (clk), .d (n_14613), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [7]));
  CDN_flop \data_stack_mem_reg[8][0] (.clk (clk), .d (n_13866), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [0]));
  CDN_flop \data_stack_mem_reg[8][1] (.clk (clk), .d (n_13864), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [1]));
  CDN_flop \data_stack_mem_reg[8][2] (.clk (clk), .d (n_13865), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [2]));
  CDN_flop \data_stack_mem_reg[8][3] (.clk (clk), .d (n_13863), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [3]));
  CDN_flop \data_stack_mem_reg[8][4] (.clk (clk), .d (n_13867), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [4]));
  CDN_flop \data_stack_mem_reg[8][5] (.clk (clk), .d (n_13861), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [5]));
  CDN_flop \data_stack_mem_reg[8][6] (.clk (clk), .d (n_13862), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [6]));
  CDN_flop \data_stack_mem_reg[8][7] (.clk (clk), .d (n_13860), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [7]));
  CDN_flop \data_stack_pointer_reg[0] (.clk (clk), .d (n_14678), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[0]));
  CDN_flop \data_stack_pointer_reg[1] (.clk (clk), .d (n_14679), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[1]));
  CDN_flop \data_stack_pointer_reg[2] (.clk (clk), .d (n_14682), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[2]));
  CDN_flop \data_stack_pointer_reg[3] (.clk (clk), .d (n_14681), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[3]));
  CDN_flop dout_valid_reg(.clk (clk), .d (n_13908), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (dout_valid));
  or g16632 (n_13868, data_stack_pointer[3], data_stack_pointer[0]);
  or g21335 (n_13926, wc, n_13925);
  not gc (wc, \data_stack_mem[3] [0]);
  or g21355 (n_13934, wc0, n_13933);
  not gc0 (wc0, \data_stack_mem[7] [0]);
  or g22075 (n_13828, enable_n, n_13827);
  nand g25466 (n_13973, n_13919, \data_stack_mem[2] [1]);
  nand g25486 (n_14103, n_13919, \data_stack_mem[2] [3]);
  nand g25492 (n_14307, n_13919, \data_stack_mem[2] [6]);
  nand g25498 (n_13966, n_13929, \data_stack_mem[5] [0]);
  nand g25502 (n_13968, n_13927, \data_stack_mem[4] [0]);
  nand g25506 (n_14376, n_13919, \data_stack_mem[2] [7]);
  nand g25512 (n_13964, n_13931, \data_stack_mem[6] [0]);
  nand g25516 (n_13970, n_13925, \data_stack_mem[3] [0]);
  nand g25523 (n_13961, n_13933, \data_stack_mem[7] [0]);
  nand g25527 (n_14011, n_13935, \data_stack_mem[8] [0]);
  or g25542 (n_14451, n_14449, n_14450);
  or g25543 (n_14506, n_14451, n_14505);
  nand g25547 (n_14173, n_13919, \data_stack_mem[2] [4]);
  nand g25553 (n_13974, n_13923, \data_stack_mem[2] [0]);
  or g25605 (n_13922, \data_stack_mem[0] [0], wc1);
  not gc1 (wc1, \data_stack_mem[1] [0]);
  or g25642 (n_14607, wc2, data_stack_pointer[3]);
  not gc2 (wc2, data_stack_pointer[0]);
  or g25670 (n_14408, wc3, n_14407);
  not gc3 (wc3, n_14402);
  or g25693 (n_14502, n_14457, n_14439);
  or g25814 (n_14454, n_14453, n_14452);
  or g25833 (n_14456, n_14440, n_14455);
  nand g25951 (n_14241, n_13919, \data_stack_mem[2] [5]);
  nand g25957 (n_14024, n_13919, \data_stack_mem[2] [2]);
  nand g26022 (n_14233, data_stack_pointer[3], \data_stack_mem[7] [5]);
  or g26060 (n_13826, sh_bit_cnt[0], sh_bit_cnt[1]);
  or g26061 (n_13827, n_13826, sh_bit_cnt[2]);
  nand g26064 (n_13962, data_stack_pointer[3], \data_stack_mem[7] [1]);
  or g26086 (n_14415, n_14409, n_14414);
  or g26088 (n_14578, wc4, n_13853);
  not gc4 (wc4, sh_reg_in[8]);
  or g26104 (n_13813, sh_reg_out_bit_counter[0],
       sh_reg_out_bit_counter[1]);
  or g26105 (n_13814, n_13813, sh_reg_out_bit_counter[2]);
  or g26108 (n_13869, n_13868, data_stack_pointer[2]);
  or g26109 (n_13870, n_13869, data_stack_pointer[1]);
  or g26113 (n_13815, n_13814, sh_reg_out_bit_counter[3]);
  or g26153 (n_14608, wc5, n_14607);
  not gc5 (wc5, data_stack_pointer[2]);
  or g26206 (n_14508, n_14507, n_14454);
  nand g26263 (n_14208, data_stack_pointer[3], \data_stack_mem[7] [4]);
  or g26271 (n_13874, n_13872, sh_reg_in[4]);
  or g26283 (n_14446, n_14444, n_14445);
  or g26291 (n_14448, n_14447, n_14441);
  or g26295 (n_14510, n_14509, n_14456);
  nand g26417 (n_13825, out_fifo_write_pointer[2],
       out_fifo_write_pointer[1]);
  or g26418 (n_13830, n_13825, n_13829);
  or g26419 (n_13833, n_13825, n_13832);
  or g26686 (n_13840, n_13839, n_13829);
  or g26687 (n_13842, n_13839, n_13832);
  or g26817 (n_14411, wc6, \data_stack_mem[7] [7]);
  not gc6 (wc6, data_stack_pointer[3]);
  or g26818 (n_14322, wc7, \data_stack_mem[7] [6]);
  not gc7 (wc7, data_stack_pointer[3]);
  or g26819 (n_14118, wc8, \data_stack_mem[7] [3]);
  not gc8 (wc8, data_stack_pointer[3]);
  or g26824 (n_13839, out_fifo_write_pointer[2], wc9);
  not gc9 (wc9, out_fifo_write_pointer[1]);
  or g26842 (n_14672, n_13851, wc10);
  not gc10 (wc10, out_fifo_read_pointer[0]);
  or g26857 (n_14178, n_13920, wc11);
  not gc11 (wc11, \data_stack_mem[0] [4]);
  or g26870 (n_14462, n_13918, wc12);
  not gc12 (wc12, \data_stack_mem[4] [7]);
  or g26874 (n_13999, n_13918, wc13);
  not gc13 (wc13, \data_stack_mem[4] [1]);
  or g26883 (n_14275, n_13918, wc14);
  not gc14 (wc14, \data_stack_mem[4] [5]);
  or g26923 (n_13924, n_13923, wc15);
  not gc15 (wc15, \data_stack_mem[2] [0]);
  or g26991 (n_13928, n_13927, wc16);
  not gc16 (wc16, \data_stack_mem[4] [0]);
  or g27028 (n_13930, n_13929, wc17);
  not gc17 (wc17, \data_stack_mem[5] [0]);
  or g27047 (n_13932, n_13931, wc18);
  not gc18 (wc18, \data_stack_mem[6] [0]);
  or g27140 (n_14494, n_14393, wc19);
  not gc19 (wc19, n_14399);
  or g27164 (n_14492, n_14391, wc20);
  not gc20 (wc20, n_14401);
  not g32605 (n_13823, rst_n);
  not g32606 (n_13824, enable_n);
  not g32607 (n_13831, n_13830);
  not g32608 (n_13834, n_13833);
  not g32609 (n_13836, n_13835);
  not g32610 (n_13838, n_13837);
  not g32611 (n_13841, n_13840);
  not g32612 (n_13843, n_13842);
  not g32613 (n_13845, n_13844);
  not g32614 (n_13847, n_13846);
  or g32622 (n_13872, sh_reg_in[0], sh_reg_in[1]);
  or g32645 (n_13936, n_13935, wc21);
  not gc21 (wc21, \data_stack_mem[8] [0]);
  or g32663 (n_13963, wc22, \data_stack_mem[7] [1]);
  not gc22 (wc22, data_stack_pointer[3]);
  or g32667 (n_13975, wc23, \data_stack_mem[2] [1]);
  not gc23 (wc23, n_13919);
  nand g32671 (n_14015, data_stack_pointer[3], \data_stack_mem[7] [2]);
  or g32672 (n_14020, n_13918, \data_stack_mem[4] [2]);
  or g32673 (n_14021, n_13918, wc24);
  not gc24 (wc24, \data_stack_mem[4] [2]);
  or g32674 (n_14025, wc25, \data_stack_mem[2] [2]);
  not gc25 (wc25, n_13919);
  or g32675 (n_14037, wc26, \data_stack_mem[7] [2]);
  not gc26 (wc26, data_stack_pointer[3]);
  nand g32691 (n_14094, data_stack_pointer[3], \data_stack_mem[7] [3]);
  or g32692 (n_14099, n_13918, \data_stack_mem[4] [3]);
  or g32693 (n_14100, n_13918, wc27);
  not gc27 (wc27, \data_stack_mem[4] [3]);
  or g32695 (n_14104, wc28, \data_stack_mem[2] [3]);
  not gc28 (wc28, n_13919);
  or g32705 (n_14169, n_13918, \data_stack_mem[4] [4]);
  or g32706 (n_14170, n_13918, wc29);
  not gc29 (wc29, \data_stack_mem[4] [4]);
  or g32708 (n_14174, wc30, \data_stack_mem[2] [4]);
  not gc30 (wc30, n_13919);
  or g32719 (n_14234, wc31, \data_stack_mem[7] [5]);
  not gc31 (wc31, data_stack_pointer[3]);
  or g32723 (n_14242, wc32, \data_stack_mem[2] [5]);
  not gc32 (wc32, n_13919);
  nand g32733 (n_14298, data_stack_pointer[3], \data_stack_mem[7] [6]);
  or g32734 (n_14303, n_13918, \data_stack_mem[4] [6]);
  or g32735 (n_14304, n_13918, wc33);
  not gc33 (wc33, \data_stack_mem[4] [6]);
  or g32737 (n_14308, wc34, \data_stack_mem[2] [6]);
  not gc34 (wc34, n_13919);
  or g32749 (n_14377, wc35, \data_stack_mem[2] [7]);
  not gc35 (wc35, n_13919);
  nand g32756 (n_14410, data_stack_pointer[3], \data_stack_mem[7] [7]);
  or g33072 (n_13940, n_13872, wc36);
  not gc36 (wc36, sh_reg_in[4]);
  or g33298 (n_14512, n_14415, wc37);
  not gc37 (wc37, n_14501);
  or g33496 (n_14883, n_13918, \data_stack_mem[4] [5]);
  or g33567 (n_14902, n_14494, wc38);
  not gc38 (wc38, n_14497);
  or g33582 (n_14909, out_fifo_write_pointer[1], wc39);
  not gc39 (wc39, out_fifo_write_pointer[2]);
  or g33583 (n_13835, n_14909, n_13829);
  or g33584 (n_13837, n_14909, n_13832);
  or g33587 (n_14910, n_14502, n_14511);
  or g33590 (n_14911, sh_reg_in[8], n_13853);
  or g33591 (n_13854, n_14911, data_stack_pointer[1]);
  or g33594 (n_14912, enable_n, n_13826);
  or g33606 (n_14916, \data_stack_mem[6] [4], n_14205);
  or g33609 (n_14917, \data_stack_mem[7] [2], n_14072);
  or g33612 (n_14918, wc40, n_14038);
  not gc40 (wc40, \data_stack_mem[7] [2]);
  or g33615 (n_14919, wc41, n_14421);
  not gc41 (wc41, \data_stack_mem[4] [7]);
  nand g33618 (n_14920, n_14370, \data_stack_mem[4] [7]);
  or g33624 (n_14922, \data_stack_mem[5] [5], n_14260);
  or g33630 (n_14924, \data_stack_mem[6] [3], n_14135);
  or g33645 (n_14929, wc42, n_14423);
  not gc42 (wc42, \data_stack_mem[3] [7]);
  nand g33651 (n_14931, \data_stack_mem[3] [7], n_14374);
  or g33657 (n_14933, wc43, n_14318);
  not gc43 (wc43, \data_stack_mem[4] [6]);
  or g33660 (n_14934, \data_stack_mem[4] [6], n_14342);
  or g33663 (n_14935, \data_stack_mem[5] [4], n_14194);
  or g33678 (n_14940, n_13932, n_13992);
  or g33681 (n_14941, n_14266, n_14267);
  or g33684 (n_14942, n_14117, n_14119);
  or g33690 (n_14944, wc44, n_14316);
  not gc44 (wc44, \data_stack_mem[3] [6]);
  or g33693 (n_14945, \data_stack_mem[3] [6], n_14343);
  or g33696 (n_14946, wc45, n_14427);
  not gc45 (wc45, \data_stack_mem[2] [7]);
  or g33702 (n_14948, \data_stack_mem[4] [4], n_14202);
  or g33708 (n_14950, \data_stack_mem[5] [2], n_14059);
  or g33714 (n_14952, wc46, n_14249);
  not gc46 (wc46, \data_stack_mem[3] [5]);
  or g33717 (n_14953, \data_stack_mem[4] [3], n_14145);
  nand g33720 (n_14954, \data_stack_mem[8] [7], n_14412);
  or g33723 (n_14955, n_14112, n_14111);
  or g33726 (n_14956, \data_stack_mem[4] [2], n_14068);
  or g33729 (n_14957, n_14261, n_14265);
  or g33732 (n_14958, n_14270, n_14271);
  nand g33738 (n_14960, \data_stack_mem[2] [7], n_14383);
  or g33741 (n_14961, wc47, n_14182);
  not gc47 (wc47, \data_stack_mem[3] [4]);
  or g33744 (n_14962, n_14512, wc48);
  not gc48 (wc48, n_14526);
  or g33753 (n_14965, wc49, n_14040);
  not gc49 (wc49, \data_stack_mem[8] [2]);
  or g33758 (n_14967, wc50, n_13918);
  not gc50 (wc50, \data_stack_mem[4] [0]);
  or g33763 (n_14969, n_14247, n_14246);
  or g33769 (n_14971, \data_stack_mem[2] [5], n_14264);
  or g33775 (n_14973, wc51, n_14419);
  not gc51 (wc51, \data_stack_mem[6] [7]);
  or g33784 (n_14976, \data_stack_mem[2] [4], n_14197);
  or g33787 (n_14977, wc52, n_14175);
  not gc52 (wc52, \data_stack_mem[2] [4]);
  or g33790 (n_14978, \data_stack_mem[3] [2], n_14061);
  or g33799 (n_14981, \data_stack_mem[2] [3], n_14142);
  or g33802 (n_14982, wc53, n_14110);
  not gc53 (wc53, \data_stack_mem[2] [3]);
  or g33808 (n_14984, \data_stack_mem[6] [2], n_14057);
  or g33811 (n_14985, \data_stack_mem[6] [5], n_14258);
  or g33814 (n_14986, wc54, n_13868);
  not gc54 (wc54, data_stack_pointer[2]);
  or g33828 (n_14991, \data_stack_mem[5] [3], n_14137);
  or g33831 (n_14992, wc55, n_14436);
  not gc55 (wc55, \data_stack_mem[7] [7]);
  nand g33834 (n_14993, n_13919, \data_stack_mem[2] [0]);
  or g33848 (n_14998, n_14408, wc56);
  not gc56 (wc56, n_14500);
  or g33851 (n_14999, n_14148, n_14149);
  or g33854 (n_15000, wc57, n_14114);
  not gc57 (wc57, \data_stack_mem[4] [3]);
  or g33867 (n_15005, n_14321, n_14323);
  or g33870 (n_15006, \data_stack_mem[2] [6], n_14344);
  nand g33873 (n_15007, n_14367, \data_stack_mem[6] [7]);
  or g33875 (n_14403, wc58, n_14970);
  not gc58 (wc58, n_15007);
  or g33888 (n_15012, wc59, n_14432);
  not gc59 (wc59, \data_stack_mem[5] [7]);
  or g33891 (n_15013, n_14352, n_14351);
  or g33900 (n_15017, n_13815, sh_reg_out_bit_counter[4]);
  or g33903 (n_13853, n_13828, sh_bit_cnt[3]);
  or g33910 (n_15020, wc60, n_14121);
  not gc60 (wc60, \data_stack_mem[8] [3]);
  nand g33916 (n_15022, data_stack_pointer[3], \data_stack_mem[7] [0]);
  or g33922 (n_15024, n_14187, n_14168);
  or g33925 (n_15025, wc61, n_14190);
  not gc61 (wc61, \data_stack_mem[8] [4]);
  or g33931 (n_15027, wc62, n_14309);
  not gc62 (wc62, \data_stack_mem[2] [6]);
  or g33934 (n_15028, \data_stack_mem[8] [6], n_14353);
  or g33937 (n_15029, wc63, n_14022);
  not gc63 (wc63, \data_stack_mem[4] [2]);
  or g33940 (n_15030, n_14492, wc64);
  not gc64 (wc64, n_14499);
  or g33946 (n_15032, \data_stack_mem[5] [6], n_14340);
  or g33951 (n_15034, \data_stack_mem[7] [4], n_14192);
  or g33954 (n_15035, \data_stack_mem[8] [2], n_14073);
  or g33960 (n_15037, \data_stack_mem[8] [5], n_14287);
  or g33963 (n_15038, out_fifo_write_pointer[1],
       out_fifo_write_pointer[2]);
  or g33964 (n_13844, n_15038, n_13829);
  or g33965 (n_13846, n_15038, n_13832);
  nand g33967 (n_15039, n_14405, \data_stack_mem[7] [7]);
  or g33976 (n_15042, \data_stack_mem[8] [3], n_14150);
  nand g33984 (n_15045, n_14368, \data_stack_mem[5] [7]);
  or g33987 (n_15046, \data_stack_mem[8] [1], wc65);
  not gc65 (wc65, n_14011);
  or g33992 (n_15048, \data_stack_mem[8] [4], n_14207);
  or g33997 (n_15050, wc66, n_13994);
  not gc66 (wc66, \data_stack_mem[8] [1]);
  or g34029 (n_14975, wc67, \data_stack_mem[0] [1]);
  not gc67 (wc67, \data_stack_mem[1] [1]);
  or g34030 (n_15009, wc68, \data_stack_mem[0] [2]);
  not gc68 (wc68, \data_stack_mem[1] [2]);
  or g34031 (n_15019, wc69, \data_stack_mem[0] [3]);
  not gc69 (wc69, \data_stack_mem[1] [3]);
  or g34032 (n_15041, wc70, \data_stack_mem[0] [4]);
  not gc70 (wc70, \data_stack_mem[1] [4]);
  or g34034 (n_14995, wc71, \data_stack_mem[0] [5]);
  not gc71 (wc71, \data_stack_mem[1] [5]);
  or g34035 (n_14989, wc72, \data_stack_mem[0] [6]);
  not gc72 (wc72, \data_stack_mem[1] [6]);
  or g34110 (n_14983, wc73, \data_stack_mem[3] [1]);
  not gc73 (wc73, n_13970);
  or g34111 (n_14930, n_13926, wc74);
  not gc74 (wc74, \data_stack_mem[3] [1]);
  or g34173 (n_15031, wc75, \data_stack_mem[4] [1]);
  not gc75 (wc75, n_13968);
  or g34174 (n_14974, n_13928, wc76);
  not gc76 (wc76, \data_stack_mem[4] [1]);
  or g34190 (n_14963, wc77, \data_stack_mem[5] [1]);
  not gc77 (wc77, n_13966);
  or g34208 (n_14943, wc78, \data_stack_mem[6] [1]);
  not gc78 (wc78, n_13964);
  or g34209 (n_14947, n_14018, wc79);
  not gc79 (wc79, \data_stack_mem[5] [2]);
  or g34232 (n_14925, wc80, \data_stack_mem[7] [1]);
  not gc80 (wc80, n_13961);
  or g34233 (n_14926, n_13934, wc81);
  not gc81 (wc81, \data_stack_mem[7] [1]);
  or g34235 (n_15023, n_14097, wc82);
  not gc82 (wc82, \data_stack_mem[5] [3]);
  or g34254 (n_14939, n_14237, wc83);
  not gc83 (wc83, \data_stack_mem[4] [5]);
  or g34262 (n_14921, n_14095, wc84);
  not gc84 (wc84, \data_stack_mem[6] [3]);
  or g34263 (n_14932, n_14186, wc85);
  not gc85 (wc85, \data_stack_mem[5] [4]);
  or g34268 (n_14496, n_14395, wc86);
  not gc86 (wc86, n_14397);
  or g34269 (n_14503, wc87, n_14443);
  not gc87 (wc87, n_14442);
  or g34297 (n_14495, n_14394, wc88);
  not gc88 (wc88, n_14398);
  or g34320 (n_15051, n_14301, wc89);
  not gc89 (wc89, \data_stack_mem[5] [6]);
  or g34322 (n_14422, n_14927, wc90);
  not gc90 (wc90, n_14919);
  or g34330 (n_15010, n_14299, wc91);
  not gc91 (wc91, \data_stack_mem[6] [6]);
  or g34335 (n_14371, n_14928, wc92);
  not gc92 (wc92, n_14920);
  or g34360 (n_14493, n_14392, wc93);
  not gc93 (wc93, n_14400);
  or g34367 (n_14420, n_15008, wc94);
  not gc94 (wc94, n_14973);
  or g34370 (n_15004, n_14493, wc95);
  not gc95 (wc95, n_14498);
  or g34556 (n_13829, n_14578, wc96);
  not gc96 (wc96, out_fifo_write_pointer[0]);
  or g34666 (n_14972, n_14139, n_14143);
  or g34679 (n_15080, n_14200, n_14196);
  or g34704 (n_15090, \data_stack_mem[6] [6], n_14339);
  or g34754 (n_14964, n_14255, n_14256);
  or g35221 (n_15313, wc97, n_14325);
  not gc97 (wc97, \data_stack_mem[8] [6]);
  or g35225 (n_15315, wc98, n_14255);
  not gc98 (wc98, \data_stack_mem[7] [5]);
  or g35227 (n_15316, wc99, n_13930);
  not gc99 (wc99, \data_stack_mem[5] [1]);
  or g35237 (n_15321, \data_stack_mem[2] [1], n_13978);
  or g35255 (n_15330, \data_stack_mem[2] [2], n_14065);
  or g35257 (n_15331, \data_stack_mem[3] [4], n_14200);
  or g35265 (n_15335, n_14232, wc100);
  not gc100 (wc100, \data_stack_mem[8] [5]);
  or g35269 (n_15337, n_14188, wc101);
  not gc101 (wc101, \data_stack_mem[7] [4]);
  or g35271 (n_15338, wc102, n_14016);
  not gc102 (wc102, \data_stack_mem[6] [2]);
  or g35275 (n_15340, wc103, n_13988);
  not gc103 (wc103, \data_stack_mem[2] [1]);
  or g35285 (n_15345, wc104, n_14183);
  not gc104 (wc104, \data_stack_mem[4] [4]);
  or g35287 (n_15346, wc105, n_14251);
  not gc105 (wc105, \data_stack_mem[5] [5]);
  or g35289 (n_15347, wc106, n_14032);
  not gc106 (wc106, \data_stack_mem[3] [2]);
  or g35321 (n_15363, wc107, n_14235);
  not gc107 (wc107, \data_stack_mem[6] [5]);
  or g35349 (n_15377, n_14031, wc108);
  not gc108 (wc108, \data_stack_mem[2] [2]);
  or g35373 (n_15389, wc109, n_14418);
  not gc109 (wc109, \data_stack_mem[8] [7]);
  or g35425 (n_15415, \data_stack_mem[0] [1], \data_stack_mem[1] [1]);
  or g35441 (n_15423, \data_stack_mem[0] [2], \data_stack_mem[1] [2]);
  or g35461 (n_15433, \data_stack_mem[0] [3], \data_stack_mem[1] [3]);
  or g35479 (n_15442, \data_stack_mem[0] [4], \data_stack_mem[1] [4]);
  or g35487 (n_15446, data_stack_pointer[1], data_stack_pointer[3]);
  or g35497 (n_15451, \data_stack_mem[0] [5], \data_stack_mem[1] [5]);
  or g35507 (n_15456, wc110, n_13937);
  not gc110 (wc110, \data_stack_mem[8] [0]);
  or g35511 (n_15458, \data_stack_mem[0] [6], \data_stack_mem[1] [6]);
  or g35535 (n_15470, sh_bit_cnt[3], n_13827);
  or g35551 (n_15478, wc111, n_13937);
  not gc111 (wc111, \data_stack_mem[8] [1]);
  or g35569 (n_15487, wc112, n_13937);
  not gc112 (wc112, \data_stack_mem[8] [5]);
  or g35573 (n_15489, \data_stack_mem[1] [1], wc113);
  not gc113 (wc113, n_13920);
  or g35575 (n_15490, \data_stack_mem[4] [1], n_13918);
  or g35577 (n_15491, \data_stack_mem[8] [1], n_13937);
  or g35601 (n_15503, \data_stack_mem[4] [7], n_13918);
  or g35605 (n_15505, \data_stack_mem[0] [0], \data_stack_mem[1] [0]);
  or g35609 (n_15507, \data_stack_mem[4] [0], n_13918);
  or g35611 (n_15508, \data_stack_mem[7] [0], wc114);
  not gc114 (wc114, data_stack_pointer[3]);
  or g35617 (n_15511, \data_stack_mem[2] [0], wc115);
  not gc115 (wc115, n_13919);
  or g35621 (n_15513, \data_stack_mem[7] [4], wc116);
  not gc116 (wc116, data_stack_pointer[3]);
  or g35625 (n_15515, \data_stack_mem[1] [5], wc117);
  not gc117 (wc117, n_13920);
  or g35627 (n_15516, \data_stack_mem[8] [5], n_13937);
  nand g39603 (n_14559, n_20744, n_20745);
  nand g39604 (n_14547, n_20708, n_20709);
  nand g39605 (n_14553, n_20726, n_20727);
  nand g39606 (n_14557, n_20738, n_20739);
  nand g39607 (n_14561, n_20750, n_20751);
  nand g39608 (n_14549, n_20714, n_20715);
  nand g39609 (n_14555, n_20732, n_20733);
  nand g39610 (n_14551, n_20720, n_20721);
  or g39611 (n_20726, n_13888, wc118);
  not gc118 (wc118, n_14546);
  or g39612 (n_20750, n_13900, wc119);
  not gc119 (wc119, n_14546);
  or g39613 (n_20744, n_13897, wc120);
  not gc120 (wc120, n_14546);
  or g39614 (n_20714, n_13882, wc121);
  not gc121 (wc121, n_14546);
  or g39615 (n_20708, n_13879, wc122);
  not gc122 (wc122, n_14546);
  or g39616 (n_20732, n_13891, wc123);
  not gc123 (wc123, n_14546);
  or g39617 (n_20720, n_13885, wc124);
  not gc124 (wc124, n_14546);
  or g39618 (n_20738, n_13894, wc125);
  not gc125 (wc125, n_14546);
  nand g39619 (n_14665, n_20762, n_20763);
  nand g39620 (n_14666, n_20768, n_20769);
  nand g39621 (n_14670, n_20792, n_20793);
  nand g39622 (n_14671, n_20798, n_20799);
  or g39623 (n_21843, wc126, n_14545);
  not gc126 (wc126, n_14542);
  or g39624 (n_21844, n_14542, wc127);
  not gc127 (wc127, n_14545);
  nand g39625 (n_14546, n_21843, n_21844);
  nand g39626 (n_14669, n_20786, n_20787);
  nand g39627 (n_14667, n_20774, n_20775);
  nand g39628 (n_14664, n_20756, n_20757);
  nand g39629 (n_14668, n_20780, n_20781);
  or g39630 (n_20780, n_13891, wc128);
  not gc128 (wc128, n_14663);
  or g39631 (n_20786, n_13894, wc129);
  not gc129 (wc129, n_14663);
  nand g39632 (n_14491, n_20432, n_20433);
  or g39633 (n_20774, n_13888, wc130);
  not gc130 (wc130, n_14663);
  or g39634 (n_20792, n_13897, wc131);
  not gc131 (wc131, n_14663);
  nand g39635 (n_14481, n_20372, n_20373);
  or g39636 (n_20768, n_13885, wc132);
  not gc132 (wc132, n_14663);
  or g39637 (n_20798, n_13900, wc133);
  not gc133 (wc133, n_14663);
  nand g39638 (n_14477, n_20348, n_20349);
  or g39639 (n_20762, n_13882, wc134);
  not gc134 (wc134, n_14663);
  nand g39640 (n_14485, n_20396, n_20397);
  nand g39641 (n_14487, n_20408, n_20409);
  or g39642 (n_20756, n_13879, wc135);
  not gc135 (wc135, n_14663);
  nand g39643 (n_14483, n_20384, n_20385);
  nand g39644 (n_14479, n_20360, n_20361);
  nand g39645 (n_14489, n_20420, n_20421);
  or g39646 (n_21845, wc136, n_14541);
  not gc136 (wc136, n_14896);
  or g39647 (n_21846, n_14896, wc137);
  not gc137 (wc137, n_14541);
  nand g39648 (n_14542, n_21845, n_21846);
  or g39649 (n_20420, n_13897, wc138);
  not gc138 (wc138, n_14476);
  or g39650 (n_21847, wc139, n_14476);
  not gc139 (wc139, n_13952);
  or g39651 (n_21848, n_13952, wc140);
  not gc140 (wc140, n_14476);
  nand g39652 (n_14541, n_21847, n_21848);
  or g39653 (n_20372, n_13885, wc141);
  not gc141 (wc141, n_14476);
  nand g39654 (n_14556, n_20690, n_20691);
  nand g39655 (n_14540, n_20660, n_20661);
  or g39656 (n_20348, n_13879, wc142);
  not gc142 (wc142, n_14476);
  nand g39657 (n_14548, n_20666, n_20667);
  or g39658 (n_20396, n_13891, wc143);
  not gc143 (wc143, n_14476);
  nand g39659 (n_14550, n_20672, n_20673);
  or g39660 (n_20384, n_13888, wc144);
  not gc144 (wc144, n_14476);
  nand g39661 (n_14552, n_20678, n_20679);
  or g39662 (n_20408, n_13894, wc145);
  not gc145 (wc145, n_14476);
  nand g39663 (n_14560, n_20702, n_20703);
  or g39664 (n_20432, n_13900, wc146);
  not gc146 (wc146, n_14476);
  or g39665 (n_20360, n_13882, wc147);
  not gc147 (wc147, n_14476);
  nand g39666 (n_14558, n_20696, n_20697);
  nand g39667 (n_21849, n_14661, n_14662);
  or g39668 (n_21850, n_14661, n_14662);
  nand g39669 (n_14663, n_21849, n_21850);
  nand g39670 (n_14554, n_20684, n_20685);
  or g39671 (n_20690, n_13894, n_14539);
  nand g39672 (n_14719, n_14715, n_20469);
  or g39673 (n_20696, n_13897, n_14539);
  or g39674 (n_20684, n_13891, n_14539);
  or g39675 (n_20702, n_13900, n_14539);
  nand g39676 (n_14721, n_14720, n_20472);
  or g39677 (n_20678, n_13888, n_14539);
  nand g39678 (n_14718, n_14715, n_20466);
  nand g39679 (n_14722, n_14720, n_20475);
  or g39680 (n_20672, n_13885, n_14539);
  nand g39681 (n_14717, n_14715, n_20463);
  nand g39682 (n_14723, n_14720, n_20478);
  or g39683 (n_20666, n_13882, n_14539);
  nand g39684 (n_14716, n_14715, n_20460);
  or g39685 (n_14476, wc148, n_20328);
  not gc148 (wc148, n_20327);
  or g39686 (n_20660, n_13879, n_14539);
  nand g39687 (n_14535, n_20645, n_20646);
  nand g39688 (n_21851, n_14458, n_14539);
  or g39689 (n_21852, n_14458, n_14539);
  nand g39690 (n_14661, n_21851, n_21852);
  nand g39691 (n_14724, n_14720, n_20481);
  nand g39692 (n_14534, n_20639, n_20640);
  nand g39693 (n_14714, n_14710, n_20457);
  nand g39694 (n_14726, n_14725, n_20484);
  nand g39695 (n_14533, n_20633, n_20634);
  nand g39696 (n_14727, n_14725, n_20487);
  nand g39697 (n_14728, n_14725, n_20490);
  nand g39698 (n_14532, n_20627, n_20628);
  nand g39699 (n_14707, n_14705, n_20439);
  nand g39700 (n_14729, n_14725, n_20493);
  nand g39701 (n_14531, n_20621, n_20622);
  nand g39702 (n_14731, n_14730, n_20496);
  nand g39703 (n_14706, n_14705, n_20436);
  nand g39704 (n_14530, n_20615, n_20616);
  nand g39705 (n_14732, n_14730, n_20499);
  nand g39706 (n_14733, n_14730, n_20502);
  nand g39707 (n_14529, n_20609, n_20610);
  nand g39708 (n_14713, n_14710, n_20454);
  nand g39709 (n_14734, n_14730, n_20505);
  nand g39710 (n_14528, n_20603, n_20604);
  nand g39711 (n_14712, n_14710, n_20451);
  nand g39712 (n_14736, n_14735, n_20508);
  nand g39713 (n_14521, n_20597, n_20598);
  nand g39714 (n_14711, n_14710, n_20448);
  nand g39715 (n_14737, n_14735, n_20511);
  nand g39716 (n_14520, n_20591, n_20592);
  nand g39717 (n_14709, n_14705, n_20445);
  nand g39718 (n_14738, n_14735, n_20514);
  nand g39719 (n_14519, n_20585, n_20586);
  nand g39720 (n_14739, n_14735, n_20517);
  nand g39721 (n_14741, n_14740, n_20520);
  nand g39722 (n_14518, n_20579, n_20580);
  nand g39723 (n_14742, n_14740, n_20523);
  nand g39724 (n_14743, n_14740, n_20526);
  nand g39725 (n_14517, n_20573, n_20574);
  nand g39726 (n_14744, n_14740, n_20529);
  nand g39727 (n_14514, n_20555, n_20556);
  nand g39728 (n_14516, n_20567, n_20568);
  nand g39729 (n_14708, n_14705, n_20442);
  nand g39730 (n_14515, n_20561, n_20562);
  nand g39731 (n_14459, n_20342, n_20343);
  or g39732 (n_20561, n_13882, n_14513);
  or g39733 (n_20567, n_13885, n_14513);
  or g39734 (n_20615, n_13885, n_14527);
  or g39735 (n_20555, n_13879, n_14513);
  or g39736 (n_20573, n_13888, n_14513);
  or g39737 (n_20639, n_13897, n_14527);
  or g39738 (n_21853, wc149, n_14527);
  not gc149 (wc149, n_14513);
  or g39739 (n_21854, n_14513, wc150);
  not gc150 (wc150, n_14527);
  nand g39740 (n_14662, n_21853, n_21854);
  or g39741 (n_14720, n_13842, n_14704);
  or g39742 (n_20579, n_13891, n_14513);
  or g39743 (n_14725, n_13830, n_14704);
  nand g39744 (n_14488, n_20414, n_20415);
  or g39745 (n_14735, n_13833, n_14704);
  or g39746 (n_20585, n_13894, n_14513);
  or g39747 (n_14740, n_13840, n_14704);
  or g39748 (n_20645, n_13900, n_14527);
  or g39749 (n_20591, n_13897, n_14513);
  or g39750 (n_14539, n_14417, n_20655);
  or g39751 (n_20597, n_13900, n_14513);
  or g39752 (n_14710, n_13835, n_14704);
  or g39753 (n_20603, n_13879, n_14527);
  nand g39754 (n_14490, n_20426, n_20427);
  or g39755 (n_20609, n_13882, n_14527);
  nand g39756 (n_14480, n_20366, n_20367);
  or g39757 (n_14705, n_13846, n_14704);
  nand g39758 (n_14478, n_20354, n_20355);
  or g39759 (n_20327, n_20324, wc151);
  not gc151 (wc151, sh_reg_in[5]);
  or g39760 (n_20621, n_13888, n_14527);
  or g39761 (n_14730, n_13844, n_14704);
  nand g39762 (n_14484, n_20390, n_20391);
  or g39763 (n_14715, n_13837, n_14704);
  or g39764 (n_20627, n_13891, n_14527);
  nand g39765 (n_14486, n_20402, n_20403);
  nand g39766 (n_14482, n_20378, n_20379);
  or g39767 (n_20633, n_13894, n_14527);
  or g39768 (n_20378, n_13888, n_14458);
  or g39769 (n_20426, n_13900, n_14458);
  or g39770 (n_14704, n_20310, wc152);
  not gc152 (wc152, rst_n);
  or g39771 (n_14527, n_14416, n_20541);
  or g39772 (n_20354, n_13882, n_14458);
  or g39773 (n_20414, n_13897, n_14458);
  or g39774 (n_20324, wc153, n_13911);
  not gc153 (wc153, n_15308);
  or g39775 (n_20402, n_13894, n_14458);
  or g39776 (n_20390, n_13891, n_14458);
  or g39777 (n_14513, n_14417, n_20550);
  or g39778 (n_20366, n_13885, n_14458);
  nand g39779 (n_20655, n_20653, n_20654);
  or g39780 (n_20342, n_13879, n_14458);
  nand g39781 (n_20550, n_20548, n_20549);
  nand g39782 (n_20654, n_15388, sh_reg_in[5]);
  or g39783 (n_20310, n_20309, wc154);
  not gc154 (wc154, sh_reg_in[5]);
  nand g39784 (n_20541, n_20539, n_20540);
  nand g39785 (n_15308, n_20300, n_20301);
  or g39786 (n_14458, n_14417, n_20337);
  or g39787 (n_20300, sh_reg_in[4], wc155);
  not gc155 (wc155, n_14460);
  or g39788 (n_20309, n_14523, n_13871);
  nand g39789 (n_20540, sh_reg_in[5], n_14523);
  nand g39790 (n_20549, n_15398, sh_reg_in[5]);
  nand g39791 (n_20337, n_20335, n_20336);
  or g39792 (n_21855, wc156, n_14910);
  not gc156 (wc156, n_14538);
  or g39793 (n_21856, n_14538, wc157);
  not gc157 (wc157, n_14910);
  nand g39794 (n_15388, n_21855, n_21856);
  or g39795 (n_20653, sh_reg_in[5], wc158);
  not gc158 (wc158, n_15387);
  nand g39796 (n_20336, n_15410, sh_reg_in[5]);
  or g39797 (n_21857, wc159, n_14289);
  not gc159 (wc159, n_14544);
  or g39798 (n_21858, n_14544, wc160);
  not gc160 (wc160, n_14289);
  nand g39799 (n_14545, n_21857, n_21858);
  nand g39800 (n_20328, n_20325, n_20326);
  or g39801 (n_21859, wc161, n_14511);
  not gc161 (wc161, n_14502);
  or g39802 (n_21860, n_14502, wc162);
  not gc162 (wc162, n_14511);
  nand g39803 (n_15398, n_21859, n_21860);
  or g39804 (n_14523, n_13874, wc163);
  not gc163 (wc163, n_20271);
  nand g39805 (n_14460, n_20255, n_20256);
  nand g39806 (n_14366, n_20249, n_20250);
  nand g39807 (n_14365, n_20243, n_20244);
  nand g39808 (n_14364, n_20237, n_20238);
  nand g39809 (n_14363, n_20231, n_20232);
  nand g39810 (n_14362, n_20225, n_20226);
  nand g39811 (n_14361, n_20219, n_20220);
  nand g39812 (n_14360, n_20213, n_20214);
  nand g39813 (n_14359, n_20207, n_20208);
  or g39814 (n_20271, n_20270, wc164);
  not gc164 (wc164, n_14439);
  or g39815 (n_20539, sh_reg_in[5], wc165);
  not gc165 (wc165, n_14962);
  or g39816 (n_20548, sh_reg_in[5], wc166);
  not gc166 (wc166, n_15397);
  nand g39817 (n_15387, n_14962, n_20532);
  or g39818 (n_21861, wc167, n_14439);
  not gc167 (wc167, n_14457);
  or g39819 (n_21862, n_14457, wc168);
  not gc168 (wc168, n_14439);
  nand g39820 (n_15410, n_21861, n_21862);
  or g39821 (n_21863, wc169, n_14155);
  not gc169 (wc169, n_14543);
  or g39822 (n_21864, n_14543, wc170);
  not gc170 (wc170, n_14155);
  nand g39823 (n_14544, n_21863, n_21864);
  or g39824 (n_20326, n_13913, wc171);
  not gc171 (wc171, n_14475);
  or g39825 (n_20255, n_13872, wc172);
  not gc172 (wc172, n_15312);
  or g39826 (n_20225, n_13888, wc173);
  not gc173 (wc173, n_14358);
  or g39827 (n_14439, n_13937, n_21024);
  or g39828 (n_20219, n_13885, wc174);
  not gc174 (wc174, n_14358);
  or g39829 (n_20249, n_13900, wc175);
  not gc175 (wc175, n_14358);
  nand g39830 (n_15397, n_14512, n_20313);
  nand g39831 (n_21865, n_15311, n_14438);
  or g39832 (n_21866, n_15311, n_14438);
  nand g39833 (n_15312, n_21865, n_21866);
  or g39834 (n_20243, n_13897, wc176);
  not gc176 (wc176, n_14358);
  or g39835 (n_20213, n_13882, wc177);
  not gc177 (wc177, n_14358);
  or g39836 (n_20335, sh_reg_in[5], wc178);
  not gc178 (wc178, n_15409);
  or g39837 (n_20237, n_13894, wc179);
  not gc179 (wc179, n_14358);
  or g39838 (n_14475, n_20294, n_20295);
  or g39839 (n_20207, n_13879, wc180);
  not gc180 (wc180, n_14358);
  or g39840 (n_20231, n_13891, wc181);
  not gc181 (wc181, n_14358);
  or g39841 (n_21867, wc182, n_14013);
  not gc182 (wc182, n_14358);
  or g39842 (n_21868, n_14358, wc183);
  not gc183 (wc183, n_14013);
  nand g39843 (n_14543, n_21867, n_21868);
  or g39844 (n_20532, wc184, n_14526);
  not gc184 (wc184, n_14512);
  or g39845 (n_14358, wc185, n_20202);
  not gc185 (wc185, n_20201);
  or g39846 (n_20313, wc186, n_14501);
  not gc186 (wc186, n_14415);
  or g39847 (n_15311, n_13937, n_20061);
  nand g39848 (n_15409, n_14415, n_20304);
  nand g39849 (n_21024, n_21023, n_20059);
  or g39850 (n_20295, wc187, n_20293);
  not gc187 (wc187, n_20292);
  or g39851 (n_20201, n_13913, wc188);
  not gc188 (wc188, n_14357);
  nand g39852 (n_14292, n_20120, n_20121);
  nand g39853 (n_20304, n_14409, n_14414);
  nand g39854 (n_14511, n_14510, n_20259);
  nand g39855 (n_14293, n_20126, n_20127);
  nand g39856 (n_20202, n_20199, n_20200);
  nand g39857 (n_14290, n_20108, n_20109);
  nand g39858 (n_20293, n_20288, n_20289);
  nand g39859 (n_14294, n_20132, n_20133);
  nand g39860 (n_14297, n_20150, n_20151);
  nand g39861 (n_14291, n_20114, n_20115);
  nand g39862 (n_21023, n_15389, n_14438);
  nand g39863 (n_21869, n_14510, n_14537);
  or g39864 (n_21870, n_14510, n_14537);
  nand g39865 (n_14538, n_21869, n_21870);
  nand g39866 (n_14295, n_20138, n_20139);
  nand g39867 (n_14296, n_20144, n_20145);
  nand g39868 (n_20061, n_15389, n_20059);
  or g39869 (n_20120, n_13885, wc189);
  not gc189 (wc189, n_14289);
  or g39870 (n_20144, n_13897, wc190);
  not gc190 (wc190, n_14289);
  or g39871 (n_20150, n_13900, wc191);
  not gc191 (wc191, n_14289);
  or g39872 (n_20059, \data_stack_mem[8] [7], wc192);
  not gc192 (wc192, n_14418);
  or g39873 (n_20114, n_13882, wc193);
  not gc193 (wc193, n_14289);
  or g39874 (n_20138, n_13894, wc194);
  not gc194 (wc194, n_14289);
  nand g39875 (n_14457, n_14456, n_20190);
  or g39876 (n_20132, n_13891, wc195);
  not gc195 (wc195, n_14289);
  or g39877 (n_20199, wc196, n_13939);
  not gc196 (wc196, n_15376);
  or g39878 (n_14414, n_13937, n_21030);
  nand g39879 (n_20259, n_14456, n_14509);
  or g39880 (n_20108, n_13879, wc197);
  not gc197 (wc197, n_14289);
  or g39881 (n_20126, n_13888, wc198);
  not gc198 (wc198, n_14289);
  or g39882 (n_14357, n_20174, n_20175);
  or g39883 (n_20288, wc199, n_14042);
  not gc199 (wc199, n_15302);
  nand g39884 (n_21030, n_21029, n_20187);
  nand g39885 (n_14438, n_20183, n_20184);
  nand g39886 (n_21871, n_14324, n_14326);
  or g39887 (n_21872, n_14324, n_14326);
  nand g39888 (n_15376, n_21871, n_21872);
  nand g39889 (n_14418, n_19915, n_21015);
  nand g39890 (n_21873, n_14413, n_14472);
  or g39891 (n_21874, n_14413, n_14472);
  nand g39892 (n_15302, n_21873, n_21874);
  or g39893 (n_14289, n_20102, n_20103);
  or g39894 (n_20270, n_20269, wc200);
  not gc200 (wc200, n_14440);
  nand g39895 (n_20190, n_14455, n_14440);
  or g39896 (n_20175, wc201, n_20173);
  not gc201 (wc201, n_20172);
  or g39897 (n_14440, n_14437, wc202);
  not gc202 (wc202, n_20067);
  nand g39901 (n_21015, n_15313, n_14324);
  or g39902 (n_20184, wc203, n_15364);
  not gc203 (wc203, n_14435);
  or g39903 (n_20183, n_14435, wc204);
  not gc204 (wc204, n_15364);
  nand g39904 (n_14472, n_14954, n_20187);
  or g39905 (n_21029, wc205, n_14413);
  not gc205 (wc205, n_14954);
  nand g39906 (n_20173, n_20168, n_20169);
  or g39907 (n_20103, n_20101, wc206);
  not gc206 (wc206, n_20100);
  or g39908 (n_14326, n_13937, n_19917);
  nand g39909 (n_19917, n_15313, n_19915);
  nand g39910 (n_20101, n_20096, n_20097);
  nand g39911 (n_21877, n_14408, n_14500);
  or g39912 (n_21878, n_14408, n_14500);
  nand g39913 (n_14501, n_21877, n_21878);
  nand g39914 (n_15364, n_19982, n_19983);
  or g39915 (n_21879, wc207, n_14506);
  not gc207 (wc207, n_14536);
  or g39916 (n_21880, n_14536, wc208);
  not gc208 (wc208, n_14506);
  nand g39917 (n_14537, n_21879, n_21880);
  or g39918 (n_20187, \data_stack_mem[8] [7], n_14412);
  or g39919 (n_20292, n_14043, wc209);
  not gc209 (wc209, n_14412);
  nand g39920 (n_14409, n_14408, n_20178);
  or g39921 (n_20168, wc210, n_14042);
  not gc210 (wc210, n_15374);
  nand g39922 (n_20067, n_14435, n_14992);
  nand g39923 (n_14437, data_stack_pointer[3], n_19986);
  or g39924 (n_14324, wc211, n_19968);
  not gc211 (wc211, n_19967);
  nand g39925 (n_14225, n_20015, n_20016);
  or g39926 (n_19983, n_14410, wc212);
  not gc212 (wc212, n_14436);
  nand g39927 (n_14509, n_14508, n_20064);
  nand g39928 (n_14230, n_20045, n_20046);
  nand g39929 (n_14224, n_20009, n_20010);
  or g39930 (n_19915, \data_stack_mem[8] [6], wc213);
  not gc213 (wc213, n_14325);
  nand g39931 (n_14231, n_20051, n_20052);
  nand g39932 (n_20102, n_20098, n_20099);
  nand g39933 (n_14412, n_20072, n_20073);
  nand g39934 (n_21881, n_14338, n_14354);
  or g39935 (n_21882, n_14338, n_14354);
  nand g39936 (n_15374, n_21881, n_21882);
  nand g39937 (n_14229, n_20039, n_20040);
  or g39938 (n_21883, wc214, n_14522);
  not gc214 (wc214, n_14508);
  or g39939 (n_21884, n_14508, wc215);
  not gc215 (wc215, n_14522);
  nand g39940 (n_14536, n_21883, n_21884);
  nand g39941 (n_14228, n_20033, n_20034);
  or g39942 (n_19982, n_14411, n_14436);
  or g39943 (n_20097, wc216, n_14914);
  not gc216 (wc216, n_15434);
  nand g39944 (n_14227, n_20027, n_20028);
  nand g39945 (n_14413, n_19977, n_21018);
  or g39946 (n_19986, \data_stack_mem[7] [7], wc217);
  not gc217 (wc217, n_14436);
  nand g39947 (n_14226, n_20021, n_20022);
  or g39948 (n_20178, n_14402, wc218);
  not gc218 (wc218, n_14407);
  nand g39949 (n_19967, n_15314, n_14321);
  nand g39950 (n_21885, n_14232, n_14273);
  or g39951 (n_21886, n_14232, n_14273);
  nand g39952 (n_15434, n_21885, n_21886);
  nand g39953 (n_14455, n_14454, n_19989);
  nand g39954 (n_14325, n_19886, n_19887);
  nand g39955 (n_20064, n_14454, n_14507);
  nand g39956 (n_14436, n_19973, n_19974);
  or g39957 (n_21887, wc219, n_14223);
  not gc219 (wc219, n_14078);
  or g39958 (n_21888, n_14078, wc220);
  not gc220 (wc220, n_14223);
  nand g39959 (n_14896, n_21887, n_21888);
  or g39960 (n_20073, wc221, n_15306);
  not gc221 (wc221, n_14404);
  or g39961 (n_14407, n_14406, wc222);
  not gc222 (wc222, n_19992);
  or g39962 (n_20051, n_13900, wc223);
  not gc223 (wc223, n_14223);
  or g39963 (n_20099, n_20094, wc224);
  not gc224 (wc224, n_13937);
  or g39964 (n_20045, n_13897, wc225);
  not gc225 (wc225, n_14223);
  or g39965 (n_20039, n_13894, wc226);
  not gc226 (wc226, n_14223);
  or g39966 (n_20033, n_13891, wc227);
  not gc227 (wc227, n_14223);
  nand g39967 (n_14354, n_15028, n_19977);
  or g39968 (n_20027, n_13888, wc228);
  not gc228 (wc228, n_14223);
  or g39969 (n_20021, n_13885, wc229);
  not gc229 (wc229, n_14223);
  nand g39970 (n_19968, n_19965, n_19966);
  or g39971 (n_20015, n_13882, wc230);
  not gc230 (wc230, n_14223);
  or g39972 (n_20072, n_14404, wc231);
  not gc231 (wc231, n_15306);
  or g39973 (n_20009, n_13879, wc232);
  not gc232 (wc232, n_14223);
  nand g39974 (n_21018, n_15028, n_14338);
  or g39978 (n_15314, n_19788, wc233);
  not gc233 (wc233, data_stack_pointer[3]);
  nand g39979 (n_19788, n_19786, n_19787);
  or g39980 (n_21891, wc234, n_14257);
  not gc234 (wc234, \data_stack_mem[8] [5]);
  or g39981 (n_21892, \data_stack_mem[8] [5], wc235);
  not gc235 (wc235, n_14257);
  nand g39982 (n_14273, n_21891, n_21892);
  nand g39983 (n_15306, n_19922, n_19923);
  or g39984 (n_20094, wc236, n_13939);
  not gc236 (wc236, n_14257);
  or g39985 (n_19965, n_14322, n_15005);
  nand g39986 (n_21893, n_14420, n_14434);
  or g39987 (n_21894, n_14420, n_14434);
  nand g39988 (n_14435, n_21893, n_21894);
  or g39989 (n_20172, n_14043, wc237);
  not gc237 (wc237, n_14353);
  nand g39990 (n_19977, \data_stack_mem[8] [6], n_14353);
  or g39991 (n_14223, wc238, n_20004);
  not gc238 (wc238, n_20003);
  or g39992 (n_19992, n_14404, wc239);
  not gc239 (wc239, n_15039);
  nand g39993 (n_19886, n_15335, n_14257);
  nand g39994 (n_14406, data_stack_pointer[3], n_19950);
  nand g39995 (n_19989, n_14453, n_14452);
  or g39996 (n_19973, \data_stack_mem[7] [6], wc240);
  not gc240 (wc240, n_15005);
  nand g39997 (n_21895, n_14492, n_14499);
  or g39998 (n_21896, n_14492, n_14499);
  nand g39999 (n_14500, n_21895, n_21896);
  or g40000 (n_20269, n_20268, wc241);
  not gc241 (wc241, n_14453);
  or g40001 (n_20096, wc242, n_14915);
  not gc242 (wc242, n_15435);
  or g40002 (n_19787, wc243, n_14323);
  not gc243 (wc243, \data_stack_mem[7] [6]);
  or g40003 (n_19786, \data_stack_mem[7] [6], wc244);
  not gc244 (wc244, n_14323);
  nand g40004 (n_14156, n_19826, n_19827);
  nand g40005 (n_14157, n_19832, n_19833);
  or g40006 (n_14257, wc245, n_19764);
  not gc245 (wc245, n_19763);
  nand g40007 (n_14158, n_19838, n_19839);
  nand g40008 (n_14159, n_19844, n_19845);
  nand g40009 (n_14160, n_19850, n_19851);
  or g40010 (n_14353, wc246, n_19902);
  not gc246 (wc246, n_19901);
  nand g40011 (n_14507, n_14506, n_19953);
  or g40012 (n_14453, n_15008, wc247);
  not gc247 (wc247, n_19875);
  nand g40013 (n_14161, n_19856, n_19857);
  or g40014 (n_19923, n_14411, wc248);
  not gc248 (wc248, n_14405);
  nand g40015 (n_14162, n_19862, n_19863);
  or g40016 (n_19966, n_19964, wc249);
  not gc249 (wc249, n_14323);
  nand g40017 (n_14163, n_19868, n_19869);
  or g40018 (n_19922, n_14410, n_14405);
  nand g40019 (n_21897, n_14391, n_14401);
  or g40020 (n_21898, n_14391, n_14401);
  nand g40021 (n_14402, n_21897, n_21898);
  nand g40022 (n_19974, n_14321, n_14323);
  nand g40023 (n_21899, n_14403, n_14390);
  or g40024 (n_21900, n_14403, n_14390);
  nand g40025 (n_14404, n_21899, n_21900);
  or g40026 (n_20003, n_13913, wc250);
  not gc250 (wc250, n_14222);
  or g40027 (n_19950, \data_stack_mem[7] [7], n_14405);
  or g40028 (n_19856, n_13894, wc251);
  not gc251 (wc251, n_14155);
  nand g40029 (n_21901, n_14272, n_14288);
  or g40030 (n_21902, n_14272, n_14288);
  nand g40031 (n_15435, n_21901, n_21902);
  nand g40034 (n_14524, n_14902, n_15004);
  or g40035 (n_19826, n_13879, wc252);
  not gc252 (wc252, n_14155);
  or g40036 (n_19862, n_13897, wc253);
  not gc253 (wc253, n_14155);
  or g40037 (n_19964, n_14321, n_14298);
  or g40038 (n_19868, n_13900, wc254);
  not gc254 (wc254, n_14155);
  nand g40039 (n_19953, n_14451, n_14505);
  nand g40040 (n_14452, n_14451, n_19872);
  nand g40041 (n_14323, n_19775, n_19776);
  nand g40042 (n_19875, n_14973, n_14434);
  nand g40043 (n_14405, n_19880, n_19881);
  or g40044 (n_14222, n_19946, n_19947);
  nand g40045 (n_19902, n_19899, n_19900);
  nand g40046 (n_19764, n_19761, n_19762);
  or g40047 (n_19832, n_13882, wc255);
  not gc255 (wc255, n_14155);
  or g40048 (n_19838, n_13885, wc256);
  not gc256 (wc256, n_14155);
  nand g40049 (n_19901, n_15375, n_14351);
  or g40050 (n_14391, n_14970, wc257);
  not gc257 (wc257, n_19800);
  or g40051 (n_15008, wc258, n_13916);
  not gc258 (wc258, n_19803);
  or g40052 (n_19844, n_13888, wc259);
  not gc259 (wc259, n_14155);
  nand g40053 (n_19763, n_15339, n_14255);
  or g40054 (n_19850, n_13891, wc260);
  not gc260 (wc260, n_14155);
  nand g40055 (n_21905, n_14300, n_14320);
  or g40056 (n_21906, n_14300, n_14320);
  nand g40057 (n_14321, n_21905, n_21906);
  or g40058 (n_15339, n_19602, wc261);
  not gc261 (wc261, data_stack_pointer[3]);
  nand g40059 (n_14338, n_19907, n_21012);
  or g40060 (n_19947, wc262, n_19945);
  not gc262 (wc262, n_19944);
  nand g40061 (n_21907, n_14493, n_14498);
  or g40062 (n_21908, n_14493, n_14498);
  nand g40063 (n_14499, n_21907, n_21908);
  or g40064 (n_14970, wc263, n_13916);
  not gc263 (wc263, n_19725);
  nand g40065 (n_14434, n_19808, n_19809);
  or g40066 (n_14155, wc264, n_19821);
  not gc264 (wc264, n_19820);
  or g40067 (n_19800, wc265, n_14390);
  not gc265 (wc265, n_15007);
  or g40068 (n_14288, n_13937, n_19908);
  or g40069 (n_19900, n_19898, wc266);
  not gc266 (wc266, n_14352);
  nand g40070 (n_19775, n_15315, n_14256);
  nand g40071 (n_20004, n_20001, n_20002);
  or g40072 (n_19899, n_14298, n_15013);
  or g40073 (n_15375, n_19797, wc267);
  not gc267 (wc267, data_stack_pointer[3]);
  or g40074 (n_19803, \data_stack_mem[6] [7], wc268);
  not gc268 (wc268, n_14419);
  or g40075 (n_20268, n_14522, wc269);
  not gc269 (wc269, n_14450);
  or g40076 (n_19762, n_19760, wc270);
  not gc270 (wc270, n_14256);
  nand g40077 (n_19872, n_14449, n_14450);
  or g40078 (n_19761, n_14234, n_14964);
  nand g40079 (n_19880, \data_stack_mem[7] [6], n_15013);
  or g40080 (n_20001, wc271, n_13939);
  not gc271 (wc271, n_15432);
  nand g40081 (n_21909, n_14392, n_14400);
  or g40082 (n_21910, n_14392, n_14400);
  nand g40083 (n_14401, n_21909, n_21910);
  nand g40084 (n_19881, n_14351, n_14352);
  or g40085 (n_19820, n_13913, wc272);
  not gc272 (wc272, n_14154);
  nand g40086 (n_14419, n_19697, n_21006);
  or g40087 (n_14450, n_14433, wc273);
  not gc273 (wc273, n_19749);
  or g40088 (n_14300, n_19698, n_13916);
  nand g40089 (n_19908, n_15037, n_19907);
  or g40090 (n_19809, wc274, n_15405);
  not gc274 (wc274, n_14431);
  or g40091 (n_19898, n_14351, n_14322);
  nand g40092 (n_19797, n_19795, n_19796);
  or g40093 (n_19808, n_14431, wc275);
  not gc275 (wc275, n_15405);
  or g40094 (n_19760, n_14255, n_14233);
  nand g40095 (n_19602, n_19600, n_19601);
  or g40096 (n_19725, \data_stack_mem[6] [7], n_14367);
  nand g40097 (n_19945, n_19940, n_19941);
  nand g40098 (n_21012, n_15037, n_14272);
  nand g40099 (n_14390, n_19730, n_19731);
  or g40100 (n_19776, \data_stack_mem[7] [5], wc276);
  not gc276 (wc276, n_14255);
  nand g40101 (n_14091, n_19679, n_19680);
  nand g40102 (n_21911, n_14189, n_14191);
  or g40103 (n_21912, n_14189, n_14191);
  nand g40104 (n_15432, n_21911, n_21912);
  nand g40105 (n_14087, n_19667, n_19668);
  nand g40106 (n_21006, n_14320, n_15010);
  or g40107 (n_14272, wc277, n_19746);
  not gc277 (wc277, n_19745);
  or g40108 (n_19600, \data_stack_mem[7] [5], wc278);
  not gc278 (wc278, n_14256);
  or g40109 (n_19601, wc279, n_14256);
  not gc279 (wc279, \data_stack_mem[7] [5]);
  nand g40110 (n_14085, n_19661, n_19662);
  nand g40111 (n_14367, n_19592, n_21000);
  nand g40112 (n_14079, n_19643, n_19644);
  or g40113 (n_19731, wc280, n_15401);
  not gc280 (wc280, n_14387);
  nand g40114 (n_15405, n_19607, n_19608);
  or g40115 (n_19795, \data_stack_mem[7] [6], n_14352);
  nand g40116 (n_19796, \data_stack_mem[7] [6], n_14352);
  nand g40117 (n_14093, n_19685, n_19686);
  or g40118 (n_19887, \data_stack_mem[8] [5], wc281);
  not gc281 (wc281, n_14232);
  nand g40119 (n_19698, n_15010, n_19697);
  nand g40120 (n_19907, \data_stack_mem[8] [5], n_14287);
  or g40121 (n_19730, n_14387, wc282);
  not gc282 (wc282, n_15401);
  nand g40122 (n_14081, n_19649, n_19650);
  or g40123 (n_19940, wc283, n_14042);
  not gc283 (wc283, n_15431);
  nand g40124 (n_19749, n_14431, n_15012);
  or g40125 (n_14154, n_19721, n_19722);
  nand g40126 (n_14083, n_19655, n_19656);
  nand g40127 (n_21913, n_15043, n_14350);
  or g40128 (n_21914, n_15043, n_14350);
  nand g40129 (n_14351, n_21913, n_21914);
  or g40130 (n_14433, wc284, n_13917);
  not gc284 (wc284, n_19620);
  or g40131 (n_14392, n_14389, wc285);
  not gc285 (wc285, n_19626);
  nand g40132 (n_14089, n_19673, n_19674);
  nand g40133 (n_14255, n_19580, n_19581);
  or g40134 (n_19581, wc286, n_15318);
  not gc286 (wc286, n_14254);
  or g40135 (n_19580, n_14254, wc287);
  not gc287 (wc287, n_15318);
  or g40136 (n_19661, n_13888, wc288);
  not gc288 (wc288, n_14078);
  nand g40137 (n_14449, n_14448, n_19623);
  or g40138 (n_19620, \data_stack_mem[5] [7], wc289);
  not gc289 (wc289, n_14432);
  nand g40139 (n_14352, n_19769, n_19770);
  or g40140 (n_15043, n_19593, n_13916);
  or g40141 (n_19655, n_13885, wc290);
  not gc290 (wc290, n_14078);
  or g40142 (n_19626, n_14387, wc291);
  not gc291 (wc291, n_15045);
  or g40143 (n_14389, wc292, n_13917);
  not gc292 (wc292, n_19572);
  or g40144 (n_19697, \data_stack_mem[6] [6], wc293);
  not gc293 (wc293, n_14299);
  or g40145 (n_19649, n_13882, wc294);
  not gc294 (wc294, n_14078);
  nand g40146 (n_14287, n_19779, n_21009);
  or g40147 (n_19685, n_13900, wc295);
  not gc295 (wc295, n_14078);
  or g40148 (n_19608, n_14369, wc296);
  not gc296 (wc296, n_14432);
  nand g40149 (n_21000, n_14350, n_15090);
  or g40150 (n_19607, n_14388, n_14432);
  or g40151 (n_19643, n_13879, wc297);
  not gc297 (wc297, n_14078);
  or g40152 (n_19667, n_13891, wc298);
  not gc298 (wc298, n_14078);
  nand g40153 (n_19745, n_15411, n_14270);
  nand g40154 (n_21915, n_14494, n_14497);
  or g40155 (n_21916, n_14494, n_14497);
  nand g40156 (n_14498, n_21915, n_21916);
  or g40157 (n_19673, n_13894, wc299);
  not gc299 (wc299, n_14078);
  nand g40158 (n_21917, n_14221, n_14218);
  or g40159 (n_21918, n_14221, n_14218);
  nand g40160 (n_15431, n_21917, n_21918);
  nand g40161 (n_19746, n_19743, n_19744);
  nand g40162 (n_14256, n_19586, n_19587);
  nand g40163 (n_14232, n_19691, n_21003);
  nand g40164 (n_21919, n_14302, n_14319);
  or g40165 (n_21920, n_14302, n_14319);
  nand g40166 (n_14320, n_21919, n_21920);
  nand g40167 (n_21921, n_14448, n_14504);
  or g40168 (n_21922, n_14448, n_14504);
  nand g40169 (n_14505, n_21921, n_21922);
  or g40170 (n_14191, n_13937, n_19692);
  or g40171 (n_19679, n_13897, wc300);
  not gc300 (wc300, n_14078);
  nand g40172 (n_15401, n_19544, n_19545);
  or g40173 (n_19722, wc301, n_19720);
  not gc301 (wc301, n_19719);
  or g40174 (n_19544, n_14369, n_14368);
  or g40175 (n_19545, n_14388, wc302);
  not gc302 (wc302, n_14368);
  or g40176 (n_19743, n_14233, n_14958);
  nand g40177 (n_21923, n_14341, n_14349);
  or g40178 (n_21924, n_14341, n_14349);
  nand g40179 (n_14350, n_21923, n_21924);
  nand g40180 (n_19946, n_19942, n_19943);
  nand g40181 (n_19821, n_19818, n_19819);
  nand g40182 (n_21925, n_14393, n_14399);
  or g40183 (n_21926, n_14393, n_14399);
  nand g40184 (n_14400, n_21925, n_21926);
  or g40185 (n_19744, n_19742, wc303);
  not gc303 (wc303, n_14271);
  nand g40186 (n_21927, n_14371, n_14386);
  or g40187 (n_21928, n_14371, n_14386);
  nand g40188 (n_14387, n_21927, n_21928);
  nand g40189 (n_21929, n_14422, n_14430);
  or g40190 (n_21930, n_14422, n_14430);
  nand g40191 (n_14431, n_21929, n_21930);
  nand g40192 (n_14432, n_19538, n_20997);
  or g40193 (n_14522, n_19575, wc304);
  not gc304 (wc304, n_14441);
  nand g40194 (n_19720, n_19715, n_19716);
  nand g40195 (n_19769, \data_stack_mem[7] [5], n_14958);
  nand g40196 (n_21009, n_15048, n_14221);
  or g40197 (n_14302, n_19539, n_13917);
  or g40198 (n_19572, \data_stack_mem[5] [7], n_14368);
  or g40199 (n_14078, wc305, n_19638);
  not gc305 (wc305, n_19637);
  nand g40200 (n_14299, n_19502, n_20985);
  nand g40201 (n_19593, n_15090, n_19592);
  or g40202 (n_15411, n_19617, wc306);
  not gc306 (wc306, data_stack_pointer[3]);
  nand g40203 (n_14218, n_15048, n_19779);
  nand g40204 (n_19623, n_14447, n_14441);
  nand g40205 (n_19692, n_15025, n_19691);
  nand g40206 (n_15318, n_19511, n_19512);
  nand g40207 (n_19586, n_15337, n_14164);
  nand g40208 (n_21003, n_14189, n_15025);
  nand g40209 (n_19592, \data_stack_mem[6] [6], n_14339);
  nand g40210 (n_19779, \data_stack_mem[8] [4], n_14207);
  or g40211 (n_14341, n_19485, n_13917);
  or g40212 (n_19818, wc307, n_13939);
  not gc307 (wc307, n_15445);
  nand g40213 (n_14368, n_19484, n_20982);
  or g40214 (n_19587, \data_stack_mem[7] [4], wc308);
  not gc308 (wc308, n_14188);
  nand g40215 (n_13960, n_19283, n_19284);
  or g40216 (n_19742, n_14270, n_14234);
  nand g40217 (n_13959, n_19277, n_19278);
  or g40218 (n_19943, wc309, n_14043);
  not gc309 (wc309, n_14207);
  or g40219 (n_19715, wc310, n_14042);
  not gc310 (wc310, n_15444);
  nand g40220 (n_13958, n_19271, n_19272);
  nand g40221 (n_13957, n_19265, n_19266);
  or g40222 (n_14393, n_14928, wc311);
  not gc311 (wc311, n_19515);
  nand g40223 (n_13956, n_19259, n_19260);
  or g40224 (n_19512, n_19510, n_13916);
  nand g40225 (n_13955, n_19253, n_19254);
  nand g40226 (n_13954, n_19247, n_19248);
  nand g40227 (n_13953, n_19241, n_19242);
  nand g40228 (n_19617, n_19615, n_19616);
  or g40229 (n_19691, \data_stack_mem[8] [4], wc312);
  not gc312 (wc312, n_14190);
  nand g40230 (n_19770, n_14270, n_14271);
  or g40231 (n_14441, n_14927, wc313);
  not gc313 (wc313, n_19518);
  nand g40232 (n_20985, n_15363, n_14254);
  or g40233 (n_19637, n_13913, wc314);
  not gc314 (wc314, n_14077);
  nand g40234 (n_20997, n_15051, n_14319);
  nand g40235 (n_19539, n_15051, n_19538);
  nand g40236 (n_21931, n_14165, n_14188);
  or g40237 (n_21932, n_14165, n_14188);
  nand g40238 (n_14189, n_21931, n_21932);
  nand g40239 (n_14221, n_19527, n_20991);
  nand g40240 (n_14339, n_19478, n_20979);
  or g40241 (n_19615, \data_stack_mem[7] [5], n_14271);
  nand g40242 (n_21933, n_14259, n_14269);
  or g40243 (n_21934, n_14259, n_14269);
  nand g40244 (n_14270, n_21933, n_21934);
  or g40245 (n_19265, n_13891, wc315);
  not gc315 (wc315, n_13952);
  or g40246 (n_19538, \data_stack_mem[5] [6], wc316);
  not gc316 (wc316, n_14301);
  nand g40247 (n_21935, n_14120, n_14122);
  or g40248 (n_21936, n_14120, n_14122);
  nand g40249 (n_15445, n_21935, n_21936);
  or g40250 (n_19271, n_13894, wc317);
  not gc317 (wc317, n_13952);
  or g40251 (n_19283, n_13900, wc318);
  not gc318 (wc318, n_13952);
  or g40252 (n_19515, wc319, n_14386);
  not gc319 (wc319, n_14920);
  or g40253 (n_14188, wc320, n_19368);
  not gc320 (wc320, n_19367);
  nand g40254 (n_21937, n_14134, n_14151);
  or g40255 (n_21938, n_14134, n_14151);
  nand g40256 (n_15444, n_21937, n_21938);
  or g40257 (n_19277, n_13897, wc321);
  not gc321 (wc321, n_13952);
  nand g40258 (n_14190, n_19523, n_20988);
  nand g40259 (n_19518, n_14919, n_14430);
  nand g40260 (n_21939, n_14193, n_14206);
  or g40261 (n_21940, n_14193, n_14206);
  nand g40262 (n_14207, n_21939, n_21940);
  or g40263 (n_19502, \data_stack_mem[6] [5], wc322);
  not gc322 (wc322, n_14235);
  nand g40264 (n_19616, \data_stack_mem[7] [5], n_14271);
  nand g40265 (n_19485, n_15032, n_19484);
  or g40266 (n_14927, n_13918, wc323);
  not gc323 (wc323, n_19299);
  or g40267 (n_14928, n_13918, wc324);
  not gc324 (wc324, n_19308);
  or g40268 (n_19241, n_13879, wc325);
  not gc325 (wc325, n_13952);
  or g40269 (n_14165, n_19494, wc326);
  not gc326 (wc326, data_stack_pointer[3]);
  or g40270 (n_14077, n_19568, n_19569);
  or g40271 (n_19247, n_13882, wc327);
  not gc327 (wc327, n_13952);
  nand g40272 (n_20982, n_15032, n_14349);
  or g40273 (n_19253, n_13885, wc328);
  not gc328 (wc328, n_13952);
  or g40274 (n_19511, n_14877, n_14235);
  or g40275 (n_19259, n_13888, wc329);
  not gc329 (wc329, n_13952);
  nand g40276 (n_19510, n_14235, \data_stack_mem[6] [5]);
  nand g40277 (n_19368, n_19365, n_19366);
  nand g40278 (n_14301, n_19373, n_19374);
  nand g40279 (n_20979, n_14985, n_14269);
  nand g40280 (n_14349, n_19319, n_19320);
  nand g40281 (n_14092, n_19472, n_19473);
  nand g40282 (n_14090, n_19466, n_19467);
  nand g40283 (n_14088, n_19460, n_19461);
  nand g40284 (n_14086, n_19454, n_19455);
  nand g40285 (n_14447, n_14446, n_19296);
  nand g40286 (n_20988, n_15020, n_14120);
  nand g40287 (n_14271, n_19532, n_20994);
  nand g40288 (n_14254, n_19211, n_19212);
  nand g40289 (n_14084, n_19448, n_19449);
  nand g40290 (n_14082, n_19442, n_19443);
  nand g40291 (n_14319, n_19346, n_19347);
  or g40292 (n_19569, wc330, n_19567);
  not gc330 (wc330, n_19566);
  nand g40293 (n_14151, n_15042, n_19527);
  nand g40294 (n_21941, n_14446, n_14503);
  or g40295 (n_21942, n_14446, n_14503);
  nand g40296 (n_14504, n_21941, n_21942);
  or g40297 (n_19308, \data_stack_mem[4] [7], n_14370);
  nand g40298 (n_14235, n_19379, n_19380);
  nand g40299 (n_19484, \data_stack_mem[5] [6], n_14340);
  or g40300 (n_13952, wc331, n_19236);
  not gc331 (wc331, n_19235);
  nand g40301 (n_19494, n_19492, n_19493);
  or g40302 (n_14122, n_13937, n_19524);
  nand g40303 (n_14014, n_19430, n_19431);
  or g40304 (n_14259, n_19479, n_13916);
  nand g40305 (n_14080, n_19436, n_19437);
  or g40306 (n_14193, n_19533, wc332);
  not gc332 (wc332, data_stack_pointer[3]);
  or g40307 (n_19299, \data_stack_mem[4] [7], wc333);
  not gc333 (wc333, n_14421);
  nand g40308 (n_20991, n_15042, n_14134);
  nand g40309 (n_19638, n_19635, n_19636);
  nand g40310 (n_19527, \data_stack_mem[8] [3], n_14150);
  nand g40311 (n_19236, n_19233, n_19234);
  or g40312 (n_14120, wc334, n_19341);
  not gc334 (wc334, n_19340);
  nand g40313 (n_20994, n_15034, n_14206);
  nand g40316 (n_14497, n_14496, n_14495);
  nand g40317 (n_19479, n_14985, n_19478);
  nand g40318 (n_19533, n_15034, n_19532);
  or g40319 (n_19365, n_14167, n_15024);
  or g40320 (n_19493, wc335, n_14164);
  not gc335 (wc335, \data_stack_mem[7] [4]);
  nand g40321 (n_14421, n_19205, n_20970);
  nand g40322 (n_14269, n_19313, n_19314);
  or g40323 (n_19379, \data_stack_mem[6] [4], wc336);
  not gc336 (wc336, n_15024);
  or g40324 (n_19635, wc337, n_13939);
  not gc337 (wc337, n_15449);
  or g40325 (n_19211, n_14251, wc338);
  not gc338 (wc338, n_15361);
  or g40326 (n_19212, wc339, n_15361);
  not gc339 (wc339, n_14251);
  nand g40327 (n_19296, n_14444, n_14445);
  nand g40328 (n_19373, n_15346, n_14253);
  nand g40329 (n_19567, n_19562, n_19563);
  or g40330 (n_19346, n_14317, wc340);
  not gc340 (wc340, n_15400);
  or g40331 (n_19347, wc341, n_15400);
  not gc341 (wc341, n_14317);
  nand g40332 (n_14340, n_19187, n_20961);
  or g40333 (n_19430, n_13879, wc342);
  not gc342 (wc342, n_14013);
  or g40334 (n_19436, n_13882, wc343);
  not gc343 (wc343, n_14013);
  or g40335 (n_19442, n_13885, wc344);
  not gc344 (wc344, n_14013);
  or g40336 (n_19448, n_13888, wc345);
  not gc345 (wc345, n_14013);
  or g40337 (n_19454, n_13891, wc346);
  not gc346 (wc346, n_14013);
  or g40338 (n_19460, n_13894, wc347);
  not gc347 (wc347, n_14013);
  or g40339 (n_19366, n_19364, wc348);
  not gc348 (wc348, n_14168);
  or g40340 (n_19466, n_13897, wc349);
  not gc349 (wc349, n_14013);
  or g40341 (n_19492, \data_stack_mem[7] [4], wc350);
  not gc350 (wc350, n_14164);
  or g40342 (n_19472, n_13900, wc351);
  not gc351 (wc351, n_14013);
  or g40343 (n_19319, n_14348, wc352);
  not gc352 (wc352, n_15383);
  or g40344 (n_19320, wc353, n_15383);
  not gc353 (wc353, n_14348);
  nand g40345 (n_14430, n_19223, n_19224);
  or g40346 (n_19719, n_14043, wc354);
  not gc354 (wc354, n_14150);
  nand g40347 (n_14370, n_19193, n_20964);
  nand g40348 (n_19524, n_15020, n_19523);
  or g40349 (n_19575, n_14503, wc355);
  not gc355 (wc355, n_14445);
  nand g40350 (n_14164, n_19304, n_19305);
  nand g40351 (n_19532, \data_stack_mem[7] [4], n_14192);
  or g40352 (n_14150, wc356, n_19395);
  not gc356 (wc356, n_19394);
  or g40353 (n_19562, wc357, n_14042);
  not gc357 (wc357, n_15448);
  or g40354 (n_19233, n_13913, wc358);
  not gc358 (wc358, n_13951);
  nand g40355 (n_19341, n_19338, n_19339);
  nand g40356 (n_19340, n_15386, n_14117);
  or g40357 (n_19523, \data_stack_mem[8] [3], wc359);
  not gc359 (wc359, n_14121);
  nand g40358 (n_21945, n_14394, n_14398);
  or g40359 (n_21946, n_14394, n_14398);
  nand g40360 (n_14399, n_21945, n_21946);
  or g40361 (n_19364, n_14187, n_14166);
  nand g40362 (n_19478, \data_stack_mem[6] [5], n_14258);
  nand g40363 (n_14386, n_19217, n_19218);
  nand g40364 (n_19367, n_15336, n_14187);
  or g40365 (n_19313, n_14268, wc360);
  not gc360 (wc360, n_15326);
  or g40366 (n_19314, wc361, n_15326);
  not gc361 (wc361, n_14268);
  nand g40367 (n_19380, n_14187, n_14168);
  nand g40368 (n_15361, n_19103, n_19104);
  or g40369 (n_14445, n_14424, wc362);
  not gc362 (wc362, n_19170);
  nand g40370 (n_20970, n_14933, n_14317);
  or g40371 (n_19374, \data_stack_mem[5] [5], wc363);
  not gc363 (wc363, n_14251);
  or g40372 (n_14013, n_19424, n_19425);
  nand g40373 (n_15400, n_19130, n_19131);
  nand g40374 (n_20961, n_14922, n_14268);
  nand g40375 (n_15383, n_19109, n_19110);
  or g40376 (n_19224, wc364, n_15424);
  not gc364 (wc364, n_14429);
  or g40377 (n_19223, n_14429, wc365);
  not gc365 (wc365, n_15424);
  nand g40378 (n_20964, n_14934, n_14348);
  nand g40379 (n_21947, n_14039, n_14041);
  or g40380 (n_21948, n_14039, n_14041);
  nand g40381 (n_15449, n_21947, n_21948);
  nand g40382 (n_21949, n_14056, n_14074);
  or g40383 (n_21950, n_14056, n_14074);
  nand g40384 (n_15448, n_21949, n_21950);
  or g40385 (n_19205, \data_stack_mem[4] [6], wc366);
  not gc366 (wc366, n_14318);
  or g40386 (n_15336, n_19089, n_13916);
  nand g40387 (n_14134, n_19293, n_20976);
  or g40388 (n_19304, \data_stack_mem[7] [3], wc367);
  not gc367 (wc367, n_14942);
  nand g40389 (n_14192, n_19352, n_19353);
  nand g40390 (n_19395, n_19392, n_19393);
  nand g40391 (n_19394, n_15414, n_14148);
  or g40392 (n_13951, n_19157, n_19158);
  or g40393 (n_19339, n_19337, wc368);
  not gc368 (wc368, n_14119);
  or g40394 (n_19338, n_14118, n_14942);
  or g40395 (n_15386, n_19125, wc369);
  not gc369 (wc369, data_stack_pointer[3]);
  nand g40396 (n_14121, n_19289, n_20973);
  nand g40397 (n_14206, n_19325, n_19326);
  or g40398 (n_14394, n_14375, wc370);
  not gc370 (wc370, n_19161);
  nand g40399 (n_21951, n_14238, n_14250);
  or g40400 (n_21952, n_14238, n_14250);
  nand g40401 (n_14251, n_21951, n_21952);
  nand g40402 (n_14258, n_19199, n_20967);
  or g40403 (n_19218, wc371, n_15421);
  not gc371 (wc371, n_14385);
  or g40404 (n_19217, n_14385, wc372);
  not gc372 (wc372, n_15421);
  or g40405 (n_14268, wc373, n_19053);
  not gc373 (wc373, n_19052);
  nand g40406 (n_14187, n_19175, n_19176);
  nand g40407 (n_15326, n_19079, n_19080);
  or g40408 (n_19103, n_14252, n_14253);
  or g40409 (n_19104, n_14236, wc374);
  not gc374 (wc374, n_14253);
  nand g40410 (n_19170, n_14929, n_14429);
  nand g40411 (n_14424, n_13914, n_19035);
  or g40412 (n_19425, n_19423, wc375);
  not gc375 (wc375, n_19422);
  or g40413 (n_19130, n_14303, n_14318);
  or g40414 (n_19131, n_14304, wc376);
  not gc376 (wc376, n_14318);
  or g40415 (n_19109, n_14304, n_14342);
  or g40416 (n_19110, n_14303, wc377);
  not gc377 (wc377, n_14342);
  nand g40417 (n_19193, \data_stack_mem[4] [6], n_14342);
  nand g40418 (n_15424, n_19010, n_19011);
  or g40419 (n_14041, n_13937, n_19290);
  or g40420 (n_19161, wc378, n_14385);
  not gc378 (wc378, n_14931);
  or g40421 (n_19393, n_19391, wc379);
  not gc379 (wc379, n_14149);
  or g40422 (n_19079, n_14236, n_14260);
  nand g40423 (n_19290, n_14965, n_19289);
  nand g40424 (n_19352, \data_stack_mem[7] [3], n_14999);
  or g40425 (n_19392, n_14094, n_14999);
  or g40426 (n_19325, n_14204, wc380);
  not gc380 (wc380, n_15385);
  or g40427 (n_19080, n_14252, wc381);
  not gc381 (wc381, n_14260);
  nand g40428 (n_19089, n_19087, n_19088);
  or g40429 (n_15414, n_19140, wc382);
  not gc382 (wc382, data_stack_pointer[3]);
  nand g40430 (n_20973, n_14965, n_14039);
  or g40431 (n_19326, wc383, n_15385);
  not gc383 (wc383, n_14204);
  or g40432 (n_19175, n_15319, n_14185);
  nand g40433 (n_19423, n_19418, n_19419);
  nand g40434 (n_14253, n_18992, n_20949);
  nand g40435 (n_14317, n_19064, n_19065);
  nand g40436 (n_20976, n_15035, n_14056);
  nand g40437 (n_14342, n_19070, n_19071);
  nand g40438 (n_15421, n_19004, n_19005);
  nand g40439 (n_14318, n_18980, n_20943);
  nand g40440 (n_19052, n_15329, n_14266);
  nand g40441 (n_19125, n_19123, n_19124);
  or g40442 (n_19010, n_14372, n_14423);
  nand g40443 (n_19176, n_14185, n_15319);
  or g40444 (n_19011, n_14373, wc384);
  not gc384 (wc384, n_14423);
  nand g40445 (n_20967, n_14204, n_14916);
  or g40446 (n_14238, n_13918, n_18981);
  or g40447 (n_19337, n_14117, n_14094);
  nand g40448 (n_14074, n_15035, n_19293);
  nand g40449 (n_19305, n_14117, n_14119);
  nand g40450 (n_19157, n_19153, n_19154);
  nand g40451 (n_19187, \data_stack_mem[5] [5], n_14260);
  nand g40452 (n_19053, n_19050, n_19051);
  nand g40453 (n_14375, n_13914, n_19032);
  or g40454 (n_19035, \data_stack_mem[3] [7], wc385);
  not gc385 (wc385, n_14423);
  or g40455 (n_19065, wc386, n_15417);
  not gc386 (wc386, n_14315);
  nand g40456 (n_21953, n_14195, n_14203);
  or g40457 (n_21954, n_14195, n_14203);
  nand g40458 (n_14204, n_21953, n_21954);
  nand g40459 (n_19140, n_19138, n_19139);
  or g40460 (n_19391, n_14148, n_14118);
  or g40461 (n_19418, wc387, n_14915);
  not gc387 (wc387, n_15453);
  or g40462 (n_19419, wc388, n_14914);
  not gc388 (wc388, n_15452);
  nand g40463 (n_19293, \data_stack_mem[8] [2], n_14073);
  nand g40464 (n_18981, n_14939, n_18980);
  or g40465 (n_15329, n_13918, n_18897);
  nand g40466 (n_14423, n_18914, n_20931);
  nand g40467 (n_19353, n_14148, n_14149);
  or g40468 (n_19050, n_19048, wc389);
  not gc389 (wc389, n_14267);
  or g40469 (n_19289, \data_stack_mem[8] [2], wc390);
  not gc390 (wc390, n_14040);
  or g40470 (n_19051, n_14941, n_14275);
  nand g40471 (n_14260, n_18974, n_20940);
  nand g40472 (n_19070, \data_stack_mem[4] [5], n_14941);
  nand g40473 (n_14348, n_19058, n_19059);
  or g40474 (n_19154, wc391, n_13942);
  not gc391 (wc391, n_15454);
  nand g40475 (n_20949, n_14932, n_14185);
  or g40476 (n_19124, wc392, n_14119);
  not gc392 (wc392, \data_stack_mem[7] [3]);
  or g40477 (n_19087, \data_stack_mem[6] [4], wc393);
  not gc393 (wc393, n_14168);
  or g40478 (n_19123, \data_stack_mem[7] [3], wc394);
  not gc394 (wc394, n_14119);
  or g40479 (n_19088, wc395, n_14168);
  not gc395 (wc395, \data_stack_mem[6] [4]);
  nand g40480 (n_14039, n_19166, n_19167);
  nand g40481 (n_15385, n_19115, n_19116);
  nand g40482 (n_21955, n_14096, n_14116);
  or g40483 (n_21956, n_14096, n_14116);
  nand g40484 (n_14117, n_21955, n_21956);
  or g40485 (n_19566, n_14043, wc396);
  not gc396 (wc396, n_14073);
  or g40486 (n_19004, n_14373, n_14374);
  or g40487 (n_19005, n_14372, wc397);
  not gc397 (wc397, n_14374);
  nand g40488 (n_20943, n_14250, n_14939);
  or g40489 (n_15319, n_18993, n_13917);
  or g40490 (n_19064, n_14315, wc398);
  not gc398 (wc398, n_15417);
  or g40491 (n_19032, \data_stack_mem[3] [7], n_14374);
  nand g40492 (n_18897, n_18895, n_18896);
  nand g40493 (n_18993, n_14932, n_18992);
  nand g40494 (n_15417, n_18848, n_18849);
  nand g40495 (n_14429, n_18944, n_18945);
  nand g40496 (n_21957, n_13936, n_13995);
  or g40497 (n_21958, n_13936, n_13995);
  nand g40498 (n_15452, n_21957, n_21958);
  nand g40499 (n_14374, n_18908, n_20928);
  nand g40500 (n_20931, n_14944, n_14315);
  or g40501 (n_19116, n_14167, wc399);
  not gc399 (wc399, n_14205);
  or g40502 (n_19167, wc400, n_15404);
  not gc400 (wc400, n_14036);
  or g40503 (n_19115, n_14166, n_14205);
  nand g40504 (n_14168, n_18986, n_20946);
  nand g40505 (n_19199, \data_stack_mem[6] [4], n_14205);
  nand g40506 (n_21959, n_14442, n_14443);
  or g40507 (n_21960, n_14442, n_14443);
  nand g40508 (n_14444, n_21959, n_21960);
  or g40509 (n_14195, n_18975, n_13917);
  or g40510 (n_19166, n_14036, wc401);
  not gc401 (wc401, n_15404);
  nand g40511 (n_21961, n_14136, n_14147);
  or g40512 (n_21962, n_14136, n_14147);
  nand g40513 (n_14148, n_21961, n_21962);
  or g40514 (n_14096, n_18987, n_13916);
  nand g40515 (n_19158, n_19155, n_19156);
  nand g40516 (n_19424, n_19420, n_19421);
  or g40517 (n_19058, n_14347, wc402);
  not gc402 (wc402, n_15413);
  nand g40518 (n_21963, n_14395, n_14397);
  or g40519 (n_21964, n_14395, n_14397);
  nand g40520 (n_14398, n_21963, n_21964);
  or g40521 (n_19059, wc403, n_15413);
  not gc403 (wc403, n_14347);
  nand g40522 (n_20940, n_14935, n_14203);
  nand g40523 (n_19071, n_14267, n_14266);
  nand g40524 (n_21965, n_13985, n_14012);
  or g40525 (n_21966, n_13985, n_14012);
  nand g40526 (n_15453, n_21965, n_21966);
  nand g40527 (n_14119, n_18998, n_20952);
  nand g40528 (n_14073, n_19181, n_19182);
  or g40529 (n_15454, wc404, n_19029);
  not gc404 (wc404, n_19028);
  nand g40530 (n_14385, n_18932, n_18933);
  nand g40531 (n_19139, \data_stack_mem[7] [3], n_14149);
  nand g40532 (n_14185, n_18866, n_18867);
  or g40533 (n_19048, n_14883, n_14266);
  or g40534 (n_19138, \data_stack_mem[7] [3], n_14149);
  nand g40535 (n_14040, n_19074, n_20958);
  or g40536 (n_18980, \data_stack_mem[4] [5], wc405);
  not gc405 (wc405, n_14237);
  or g40537 (n_18992, \data_stack_mem[5] [4], wc406);
  not gc406 (wc406, n_14186);
  or g40538 (n_18849, n_14306, wc407);
  not gc407 (wc407, n_14316);
  or g40539 (n_18848, n_14305, n_14316);
  nand g40540 (n_20928, n_14945, n_14347);
  or g40541 (n_14442, n_14428, wc408);
  not gc408 (wc408, n_18861);
  nand g40542 (n_20946, n_14116, n_14921);
  nand g40543 (n_14056, n_18962, n_20934);
  nand g40544 (n_14205, n_18968, n_20937);
  nand g40545 (n_15404, n_18902, n_18903);
  nand g40546 (n_15413, n_18842, n_18843);
  nand g40547 (n_18987, n_14921, n_18986);
  nand g40548 (n_14237, n_18878, n_18879);
  nand g40549 (n_14149, n_19016, n_20955);
  nand g40550 (n_20952, n_14036, n_14918);
  or g40551 (n_18933, n_15436, wc409);
  not gc409 (wc409, n_14382);
  or g40552 (n_18867, wc410, n_15359);
  not gc410 (wc410, n_14183);
  or g40553 (n_14266, wc411, n_18801);
  not gc411 (wc411, n_18800);
  or g40554 (n_18932, wc412, n_14382);
  not gc412 (wc412, n_15436);
  nand g40555 (n_18975, n_14935, n_18974);
  nand g40556 (n_18895, \data_stack_mem[4] [5], n_14267);
  or g40557 (n_14395, n_14384, wc413);
  not gc413 (wc413, n_18858);
  or g40558 (n_19235, n_13939, wc414);
  not gc414 (wc414, n_13938);
  nand g40559 (n_14250, n_18872, n_18873);
  or g40560 (n_18914, \data_stack_mem[3] [6], wc415);
  not gc415 (wc415, n_14316);
  or g40561 (n_19182, wc416, n_15427);
  not gc416 (wc416, n_14071);
  or g40562 (n_19181, n_14071, wc417);
  not gc417 (wc417, n_15427);
  or g40563 (n_19156, n_13940, wc418);
  not gc418 (wc418, n_13938);
  nand g40564 (n_13995, n_15050, n_19074);
  or g40565 (n_18866, n_14183, wc419);
  not gc419 (wc419, n_15359);
  or g40566 (n_14136, n_18969, n_13916);
  nand g40567 (n_19028, sh_reg_in[0], n_13938);
  or g40568 (n_18945, n_15440, wc420);
  not gc420 (wc420, n_14426);
  or g40569 (n_14012, n_13937, n_18963);
  or g40570 (n_18944, wc421, n_14426);
  not gc421 (wc421, n_15440);
  or g40571 (n_19421, n_19416, wc422);
  not gc422 (wc422, n_13937);
  nand g40572 (n_20958, n_13936, n_15050);
  nand g40573 (n_14203, n_18926, n_18927);
  or g40574 (n_18896, \data_stack_mem[4] [5], n_14267);
  nand g40575 (n_18974, \data_stack_mem[5] [4], n_14194);
  or g40576 (n_19074, \data_stack_mem[8] [1], wc423);
  not gc423 (wc423, n_13994);
  or g40577 (n_19416, wc424, n_13939);
  not gc424 (wc424, n_13994);
  nand g40578 (n_18963, n_15046, n_18962);
  or g40579 (n_18872, n_14248, wc425);
  not gc425 (wc425, n_15394);
  nand g40580 (n_14384, n_13919, n_18747);
  or g40581 (n_18858, wc426, n_14382);
  not gc426 (wc426, n_14960);
  nand g40582 (n_15427, n_18920, n_18921);
  or g40583 (n_18873, wc427, n_15394);
  not gc427 (wc427, n_14248);
  nand g40584 (n_13938, n_18950, n_18951);
  nand g40585 (n_14267, n_18830, n_20919);
  nand g40586 (n_18800, n_15334, n_14265);
  or g40587 (n_18998, \data_stack_mem[7] [2], wc428);
  not gc428 (wc428, n_14038);
  nand g40588 (n_20955, n_14071, n_14917);
  nand g40589 (n_18878, n_15345, n_14184);
  nand g40590 (n_15440, n_18743, n_18744);
  or g40591 (n_18902, n_14037, n_14038);
  or g40592 (n_18903, n_14015, wc429);
  not gc429 (wc429, n_14038);
  or g40593 (n_18986, \data_stack_mem[6] [3], wc430);
  not gc430 (wc430, n_14095);
  nand g40594 (n_20934, n_15046, n_13985);
  nand g40595 (n_18861, n_14426, n_14946);
  nand g40596 (n_14428, n_13919, n_18750);
  nand g40597 (n_14316, n_18725, n_20907);
  nand g40598 (n_14186, n_18824, n_20916);
  nand g40599 (n_18908, \data_stack_mem[3] [6], n_14343);
  nand g40600 (n_21967, n_14017, n_14035);
  or g40601 (n_21968, n_14017, n_14035);
  nand g40602 (n_14036, n_21967, n_21968);
  or g40603 (n_18842, n_14306, n_14343);
  nand g40604 (n_20937, n_14147, n_14924);
  nand g40605 (n_18969, n_14924, n_18968);
  or g40606 (n_18843, n_14305, wc431);
  not gc431 (wc431, n_14343);
  nand g40607 (n_15359, n_18713, n_18714);
  or g40608 (n_18926, n_14201, wc432);
  not gc432 (wc432, n_15328);
  or g40609 (n_18927, wc433, n_15328);
  not gc433 (wc433, n_14201);
  nand g40610 (n_15436, n_18731, n_18732);
  or g40611 (n_18920, n_14015, n_14072);
  nand g40612 (n_21969, n_14098, n_14115);
  or g40613 (n_21970, n_14098, n_14115);
  nand g40614 (n_14116, n_21969, n_21970);
  or g40615 (n_18921, n_14037, wc434);
  not gc434 (wc434, n_14072);
  or g40616 (n_18747, \data_stack_mem[2] [7], n_14383);
  nand g40617 (n_21971, n_14138, n_14146);
  or g40618 (n_21972, n_14138, n_14146);
  nand g40619 (n_14147, n_21971, n_21972);
  or g40620 (n_18962, wc435, n_14011);
  not gc435 (wc435, \data_stack_mem[8] [1]);
  nand g40621 (n_21973, n_14058, n_14070);
  or g40622 (n_21974, n_14058, n_14070);
  nand g40623 (n_14071, n_21973, n_21974);
  nand g40624 (n_18801, n_18798, n_18799);
  nand g40625 (n_14347, n_18773, n_18774);
  nand g40626 (n_13985, n_18938, n_18939);
  or g40627 (n_18743, n_14377, n_14427);
  or g40628 (n_18744, n_14376, wc436);
  not gc436 (wc436, n_14427);
  or g40629 (n_18713, n_14169, n_14184);
  nand g40630 (n_14038, n_18836, n_20922);
  nand g40631 (n_15328, n_18698, n_18699);
  nand g40632 (n_13994, n_18956, n_18957);
  nand g40633 (n_20907, n_14952, n_14248);
  nand g40634 (n_20919, n_14948, n_14201);
  or g40635 (n_18951, n_13936, n_13937);
  nand g40636 (n_19016, \data_stack_mem[7] [2], n_14072);
  or g40637 (n_18879, \data_stack_mem[4] [4], wc437);
  not gc437 (wc437, n_14183);
  or g40638 (n_14017, n_18693, n_13916);
  nand g40639 (n_14343, n_18806, n_18807);
  or g40640 (n_18750, \data_stack_mem[2] [7], wc438);
  not gc438 (wc438, n_14427);
  or g40641 (n_18731, n_14376, n_14383);
  or g40642 (n_18714, n_14170, wc439);
  not gc439 (wc439, n_14184);
  nand g40643 (n_20916, n_14115, n_15023);
  or g40644 (n_18732, n_14377, wc440);
  not gc440 (wc440, n_14383);
  nand g40645 (n_14095, n_18691, n_20904);
  nand g40646 (n_18968, \data_stack_mem[6] [3], n_14135);
  nand g40647 (n_14315, n_18779, n_18780);
  nand g40648 (n_14194, n_18818, n_20913);
  or g40649 (n_15334, wc441, n_18612);
  not gc441 (wc441, n_13914);
  nand g40650 (n_15394, n_18623, n_18624);
  nand g40651 (n_14184, n_18617, n_20892);
  nand g40652 (n_18612, n_18610, n_18611);
  nand g40653 (n_14115, n_18761, n_18762);
  or g40654 (n_18799, n_18797, wc442);
  not gc442 (wc442, n_14261);
  or g40655 (n_18773, wc443, n_14346);
  not gc443 (wc443, n_15420);
  nand g40656 (n_20922, n_13993, n_14926);
  or g40657 (n_18774, n_15420, wc444);
  not gc444 (wc444, n_14346);
  or g40658 (n_18623, n_14239, n_14249);
  nand g40659 (n_20913, n_14991, n_14146);
  or g40660 (n_18624, n_14240, wc445);
  not gc445 (wc445, n_14249);
  or g40661 (n_18698, n_14170, n_14202);
  or g40662 (n_14058, n_18813, n_13916);
  or g40663 (n_18699, n_14169, wc446);
  not gc446 (wc446, n_14202);
  nand g40664 (n_14183, n_18683, n_18684);
  nand g40665 (n_14383, n_18635, n_20898);
  nand g40666 (n_18806, \data_stack_mem[3] [5], n_14957);
  nand g40667 (n_14072, n_18854, n_20925);
  nand g40668 (n_14427, n_18641, n_20901);
  or g40669 (n_14138, n_18819, n_13917);
  or g40670 (n_14098, n_18825, n_13917);
  nand g40671 (n_18693, n_15338, n_18691);
  nand g40672 (n_18830, \data_stack_mem[4] [4], n_14202);
  or g40673 (n_14201, wc447, n_18657);
  not gc447 (wc447, n_18656);
  nand g40674 (n_18950, n_15456, n_13935);
  or g40675 (n_18957, wc448, n_15391);
  not gc448 (wc448, n_13993);
  or g40676 (n_18956, n_13993, wc449);
  not gc449 (wc449, n_15391);
  or g40677 (n_18938, wc450, n_13984);
  not gc450 (wc450, n_15439);
  or g40678 (n_18779, wc451, n_14314);
  not gc451 (wc451, n_15429);
  or g40679 (n_18780, n_15429, wc452);
  not gc452 (wc452, n_14314);
  or g40680 (n_18939, n_15439, wc453);
  not gc453 (wc453, n_13984);
  nand g40681 (n_20904, n_15338, n_14035);
  or g40682 (n_18725, \data_stack_mem[3] [5], wc454);
  not gc454 (wc454, n_14249);
  nand g40683 (n_14135, n_18812, n_20910);
  or g40684 (n_18798, n_14240, n_14957);
  nand g40685 (n_14249, n_18512, n_20880);
  nand g40686 (n_15420, n_18548, n_18549);
  nand g40687 (n_20892, n_15000, n_14113);
  or g40688 (n_18762, wc455, n_15349);
  not gc455 (wc455, n_14113);
  nand g40689 (n_13935, n_18785, n_18786);
  nand g40690 (n_15391, n_18719, n_18720);
  nand g40691 (n_14202, n_18602, n_20889);
  or g40692 (n_18684, wc456, n_15344);
  not gc456 (wc456, n_14181);
  nand g40693 (n_18807, n_14265, n_14261);
  nand g40694 (n_20898, n_15006, n_14346);
  nand g40695 (n_18825, n_15023, n_18824);
  or g40696 (n_18761, n_14113, wc457);
  not gc457 (wc457, n_15349);
  nand g40697 (n_15439, n_18737, n_18738);
  nand g40698 (n_18819, n_14991, n_18818);
  nand g40699 (n_20925, n_13984, n_14925);
  or g40700 (n_18683, n_14181, wc458);
  not gc458 (wc458, n_15344);
  or g40701 (n_18691, \data_stack_mem[6] [2], wc459);
  not gc459 (wc459, n_14016);
  or g40702 (n_18610, \data_stack_mem[3] [5], n_14261);
  or g40703 (n_14248, wc460, n_18489);
  not gc460 (wc460, n_18488);
  nand g40704 (n_14146, n_18755, n_18756);
  nand g40705 (n_18611, \data_stack_mem[3] [5], n_14261);
  nand g40706 (n_18813, n_14984, n_18812);
  or g40707 (n_13993, wc461, n_18672);
  not gc461 (wc461, n_18671);
  or g40708 (n_18797, n_14265, n_14239);
  nand g40709 (n_20901, n_15027, n_14314);
  nand g40710 (n_15429, n_18554, n_18555);
  nand g40711 (n_18656, n_15366, n_14200);
  nand g40712 (n_20910, n_14070, n_14984);
  nand g40713 (n_18488, n_15418, n_14246);
  nand g40714 (n_14261, n_18584, n_18585);
  or g40715 (n_18836, \data_stack_mem[7] [1], wc462);
  not gc462 (wc462, n_13934);
  or g40716 (n_18549, n_14308, wc463);
  not gc463 (wc463, n_14344);
  nand g40717 (n_20889, n_14953, n_14144);
  or g40718 (n_18548, n_14307, n_14344);
  nand g40719 (n_18672, n_18669, n_18670);
  nand g40720 (n_18812, \data_stack_mem[6] [2], n_14057);
  or g40721 (n_18641, \data_stack_mem[2] [6], wc464);
  not gc464 (wc464, n_14309);
  or g40722 (n_18854, wc465, n_13961);
  not gc465 (wc465, \data_stack_mem[7] [1]);
  nand g40723 (n_18671, n_15392, n_13992);
  or g40724 (n_18555, n_14307, wc466);
  not gc466 (wc466, n_14309);
  nand g40725 (n_18818, \data_stack_mem[5] [3], n_14137);
  or g40726 (n_18786, wc467, n_13934);
  not gc467 (wc467, data_stack_pointer[3]);
  or g40727 (n_18554, n_14308, n_14309);
  or g40728 (n_18719, n_13934, n_13963);
  nand g40729 (n_18657, n_18654, n_18655);
  or g40730 (n_14113, wc468, n_18405);
  not gc468 (wc468, n_18404);
  or g40731 (n_18756, wc469, n_15304);
  not gc469 (wc469, n_14144);
  nand g40732 (n_13984, n_18767, n_18768);
  nand g40733 (n_20880, n_14961, n_14181);
  nand g40734 (n_14016, n_18677, n_18678);
  or g40735 (n_18720, wc470, n_13962);
  not gc470 (wc470, n_13934);
  nand g40736 (n_15344, n_18440, n_18441);
  nand g40737 (n_21975, n_14060, n_14069);
  or g40738 (n_21976, n_14060, n_14069);
  nand g40739 (n_14070, n_21975, n_21976);
  or g40740 (n_18738, wc471, n_13962);
  not gc471 (wc471, n_13961);
  nand g40741 (n_18635, \data_stack_mem[2] [6], n_14344);
  or g40742 (n_18737, n_13961, n_13963);
  or g40743 (n_18755, n_14144, wc472);
  not gc472 (wc472, n_15304);
  nand g40744 (n_14265, n_18578, n_18579);
  or g40745 (n_15366, wc473, n_18528);
  not gc473 (wc473, n_13914);
  nand g40746 (n_21977, n_14019, n_14034);
  or g40747 (n_21978, n_14019, n_14034);
  nand g40748 (n_14035, n_21977, n_21978);
  or g40749 (n_18824, \data_stack_mem[5] [3], wc474);
  not gc474 (wc474, n_14097);
  or g40750 (n_15418, n_18360, wc475);
  not gc475 (wc475, n_13919);
  or g40751 (n_14019, n_18597, n_13917);
  nand g40752 (n_14344, n_18458, n_20877);
  nand g40753 (n_14057, n_18629, n_20895);
  or g40754 (n_14060, n_18591, n_13917);
  or g40755 (n_18767, n_13982, wc476);
  not gc476 (wc476, n_15396);
  nand g40756 (n_14137, n_18590, n_20883);
  nand g40757 (n_14309, n_18494, n_18495);
  or g40758 (n_18655, n_18653, wc477);
  not gc477 (wc477, n_14196);
  or g40759 (n_18768, wc478, n_15396);
  not gc478 (wc478, n_13982);
  or g40760 (n_18654, n_14172, n_15080);
  or g40761 (n_18677, \data_stack_mem[6] [1], wc479);
  not gc479 (wc479, n_14940);
  nand g40762 (n_14097, n_18596, n_20886);
  or g40763 (n_14144, wc480, n_18474);
  not gc480 (wc480, n_18473);
  or g40764 (n_18579, n_15381, wc481);
  not gc481 (wc481, n_14263);
  or g40765 (n_18578, wc482, n_14263);
  not gc482 (wc482, n_15381);
  nand g40766 (n_18584, n_15331, n_14196);
  or g40767 (n_18670, n_13983, n_14940);
  nand g40768 (n_18785, n_15022, n_13933);
  or g40769 (n_18669, n_18668, wc483);
  not gc483 (wc483, n_13932);
  or g40770 (n_18440, n_14171, n_14182);
  or g40771 (n_18512, \data_stack_mem[3] [4], wc484);
  not gc484 (wc484, n_14182);
  nand g40772 (n_18528, n_18526, n_18527);
  or g40773 (n_15392, n_18537, n_13916);
  nand g40774 (n_18404, n_15362, n_14111);
  nand g40775 (n_18489, n_18486, n_18487);
  or g40776 (n_18441, n_14172, wc485);
  not gc485 (wc485, n_14182);
  nand g40777 (n_18527, \data_stack_mem[3] [4], n_14196);
  nand g40778 (n_15381, n_18350, n_18351);
  nand g40779 (n_15304, n_18506, n_18507);
  or g40780 (n_18494, \data_stack_mem[2] [5], wc486);
  not gc486 (wc486, n_14969);
  nand g40781 (n_18591, n_14950, n_18590);
  or g40782 (n_18486, n_14242, n_14969);
  or g40783 (n_18668, n_13992, n_13965);
  nand g40784 (n_20895, n_13982, n_14943);
  nand g40785 (n_18597, n_14947, n_18596);
  nand g40786 (n_18405, n_18402, n_18403);
  nand g40787 (n_18360, n_18358, n_18359);
  nand g40788 (n_20883, n_14950, n_14069);
  nand g40789 (n_20877, n_14971, n_14263);
  nand g40790 (n_18473, n_15324, n_14143);
  nand g40791 (n_18537, n_18535, n_18536);
  nand g40792 (n_13933, n_18572, n_18573);
  nand g40793 (n_18585, \data_stack_mem[3] [4], n_14200);
  nand g40794 (n_15349, n_18518, n_18519);
  nand g40795 (n_14182, n_18422, n_18423);
  nand g40796 (n_20886, n_14034, n_14947);
  or g40797 (n_18526, \data_stack_mem[3] [4], n_14196);
  or g40798 (n_15362, wc487, n_18216);
  not gc487 (wc487, n_13914);
  nand g40799 (n_18678, n_13932, n_13992);
  nand g40800 (n_15396, n_18542, n_18543);
  or g40801 (n_18653, n_14171, n_14200);
  or g40802 (n_18422, \data_stack_mem[3] [3], wc488);
  not gc488 (wc488, n_14955);
  or g40803 (n_18402, n_14101, n_14955);
  nand g40804 (n_14181, n_18410, n_18411);
  nand g40805 (n_14034, n_18560, n_18561);
  or g40806 (n_18596, \data_stack_mem[5] [2], wc489);
  not gc489 (wc489, n_14018);
  or g40807 (n_18487, n_18485, wc490);
  not gc490 (wc490, n_14247);
  or g40808 (n_15324, wc491, n_18333);
  not gc491 (wc491, n_13914);
  or g40809 (n_18535, \data_stack_mem[6] [1], wc492);
  not gc492 (wc492, n_13932);
  or g40810 (n_18536, wc493, n_13932);
  not gc493 (wc493, \data_stack_mem[6] [1]);
  or g40811 (n_18359, wc494, n_14247);
  not gc494 (wc494, \data_stack_mem[2] [5]);
  or g40812 (n_18358, \data_stack_mem[2] [5], wc495);
  not gc495 (wc495, n_14247);
  nand g40813 (n_18458, \data_stack_mem[2] [5], n_14264);
  or g40814 (n_18629, wc496, n_13964);
  not gc496 (wc496, \data_stack_mem[6] [1]);
  nand g40815 (n_14196, n_18500, n_18501);
  nand g40816 (n_18216, n_18214, n_18215);
  or g40817 (n_18617, \data_stack_mem[4] [3], wc497);
  not gc497 (wc497, n_14114);
  nand g40818 (n_18590, \data_stack_mem[5] [2], n_14059);
  or g40819 (n_18507, n_14099, wc498);
  not gc498 (wc498, n_14145);
  or g40820 (n_18506, n_14100, n_14145);
  or g40821 (n_18542, n_13964, n_13983);
  or g40822 (n_18543, wc499, n_13965);
  not gc499 (wc499, n_13964);
  nand g40823 (n_18602, \data_stack_mem[4] [3], n_14145);
  nand g40824 (n_18495, n_14246, n_14247);
  nand g40825 (n_21979, n_13986, n_13991);
  or g40826 (n_21980, n_13986, n_13991);
  nand g40827 (n_13992, n_21979, n_21980);
  or g40828 (n_18573, n_13932, n_13916);
  nand g40829 (n_21981, n_13967, n_13981);
  or g40830 (n_21982, n_13967, n_13981);
  nand g40831 (n_13982, n_21981, n_21982);
  nand g40832 (n_14200, n_18428, n_18429);
  or g40833 (n_20100, sh_reg_in[4], n_20095);
  nand g40834 (n_14069, n_18566, n_18567);
  nand g40835 (n_18474, n_18471, n_18472);
  or g40836 (n_18350, n_14241, n_14264);
  or g40837 (n_18351, n_14242, wc500);
  not gc500 (wc500, n_14264);
  or g40838 (n_18519, n_14100, wc501);
  not gc501 (wc501, n_14114);
  or g40839 (n_18518, n_14099, n_14114);
  nand g40840 (n_14059, n_18434, n_20868);
  nand g40841 (n_14114, n_18446, n_20871);
  nand g40842 (n_18572, n_14937, n_13931);
  or g40843 (n_18403, n_18401, wc502);
  not gc502 (wc502, n_14112);
  or g40844 (n_18428, n_14199, wc503);
  not gc503 (wc503, n_15333);
  or g40845 (n_18410, n_14180, wc504);
  not gc504 (wc504, n_15408);
  nand g40846 (n_14264, n_18206, n_20859);
  or g40847 (n_18567, wc505, n_15355);
  not gc505 (wc505, n_14067);
  or g40848 (n_18566, n_14067, wc506);
  not gc506 (wc506, n_15355);
  nand g40849 (n_18500, \data_stack_mem[3] [3], n_14972);
  or g40850 (n_18429, wc507, n_15333);
  not gc507 (wc507, n_14199);
  or g40851 (n_18214, \data_stack_mem[3] [3], wc508);
  not gc508 (wc508, n_14112);
  or g40852 (n_20095, wc509, n_13913);
  not gc509 (wc509, n_14286);
  or g40853 (n_18561, wc510, n_15353);
  not gc510 (wc510, n_14033);
  or g40854 (n_13986, n_18324, n_13917);
  or g40855 (n_18215, wc511, n_14112);
  not gc511 (wc511, \data_stack_mem[3] [3]);
  or g40856 (n_18472, n_18470, wc512);
  not gc512 (wc512, n_14139);
  nand g40857 (n_14247, n_18221, n_20862);
  or g40858 (n_14382, wc513, n_16398);
  not gc513 (wc513, n_14381);
  or g40859 (n_18471, n_14102, n_14972);
  or g40860 (n_13967, n_18435, n_13917);
  or g40861 (n_18411, wc514, n_15408);
  not gc514 (wc514, n_14180);
  or g40862 (n_19422, sh_reg_in[4], n_19417);
  nand g40863 (n_18333, n_18331, n_18332);
  nand g40864 (n_18423, n_14111, n_14112);
  nand g40865 (n_14018, n_18322, n_20865);
  or g40866 (n_18560, n_14033, wc515);
  not gc515 (wc515, n_15353);
  or g40867 (n_14426, wc516, n_16410);
  not gc516 (wc516, n_14381);
  nand g40868 (n_14145, n_18452, n_20874);
  or g40869 (n_18401, n_14111, n_14102);
  nand g40870 (n_15333, n_18122, n_18123);
  nand g40871 (n_19721, n_19717, n_19718);
  nand g40872 (n_15355, n_18344, n_18345);
  or g40873 (n_14286, wc517, n_18390);
  not gc517 (wc517, n_18389);
  nand g40874 (n_20859, n_14976, n_14199);
  nand g40875 (n_18324, n_15316, n_18322);
  or g40876 (n_18470, n_14143, n_14101);
  nand g40877 (n_20174, n_20170, n_20171);
  or g40878 (n_19417, wc518, n_13913);
  not gc518 (wc518, n_14010);
  nand g40879 (n_20874, n_14067, n_14956);
  nand g40880 (n_20865, n_15316, n_13991);
  nand g40881 (n_14112, n_18182, n_18183);
  nand g40882 (n_13931, n_18416, n_18417);
  nand g40883 (n_20868, n_13981, n_14963);
  nand g40884 (n_20862, n_14977, n_14180);
  nand g40885 (n_20294, n_20290, n_20291);
  or g40886 (n_18331, \data_stack_mem[3] [3], n_14139);
  nand g40887 (n_18332, \data_stack_mem[3] [3], n_14139);
  nand g40888 (n_18435, n_14963, n_18434);
  nand g40889 (n_19568, n_19564, n_19565);
  nand g40890 (n_16410, n_16408, n_16409);
  nand g40891 (n_15353, n_18338, n_18339);
  nand g40892 (n_15408, n_18146, n_18147);
  nand g40893 (n_16398, n_16396, n_16397);
  nand g40894 (n_18501, n_14143, n_14139);
  nand g40895 (n_20871, n_15029, n_14033);
  or g40896 (n_14346, wc519, n_16314);
  not gc519 (wc519, n_14312);
  or g40897 (n_18339, n_14021, wc520);
  not gc520 (wc520, n_14022);
  or g40898 (n_18338, n_14020, n_14022);
  nand g40899 (n_21983, n_13969, n_13980);
  or g40900 (n_21984, n_13969, n_13980);
  nand g40901 (n_13981, n_21983, n_21984);
  nand g40902 (n_14033, n_18314, n_18315);
  or g40903 (n_20291, n_13942, wc521);
  not gc521 (wc521, n_14471);
  nand g40904 (n_18182, n_15347, n_14023);
  nand g40905 (n_18452, \data_stack_mem[4] [2], n_14068);
  or g40906 (n_18147, n_14173, wc522);
  not gc522 (wc522, n_14175);
  or g40907 (n_18146, n_14174, n_14175);
  or g40908 (n_18122, n_14173, n_14197);
  or g40909 (n_19565, n_13942, wc523);
  not gc523 (wc523, n_14055);
  or g40910 (n_18123, n_14174, wc524);
  not gc524 (wc524, n_14197);
  or g40911 (n_18434, wc525, n_13966);
  not gc525 (wc525, \data_stack_mem[5] [1]);
  or g40912 (n_19944, n_13942, wc526);
  not gc526 (wc526, n_14217);
  or g40913 (n_14314, wc527, n_16302);
  not gc527 (wc527, n_14312);
  or g40914 (n_14010, wc528, n_18375);
  not gc528 (wc528, n_18374);
  or g40915 (n_16409, n_16407, wc529);
  not gc529 (wc529, n_13920);
  or g40916 (n_18417, n_13930, n_13917);
  nand g40917 (n_14111, n_18176, n_18177);
  nand g40918 (n_14143, n_18170, n_18171);
  nand g40919 (n_14443, n_16421, n_16422);
  nand g40920 (n_21985, n_14062, n_14066);
  or g40921 (n_21986, n_14062, n_14066);
  nand g40922 (n_14067, n_21985, n_21986);
  or g40923 (n_18221, \data_stack_mem[2] [4], wc530);
  not gc530 (wc530, n_14175);
  nand g40924 (n_18390, n_18387, n_18388);
  or g40925 (n_18344, n_14021, n_14068);
  or g40926 (n_18345, n_14020, wc531);
  not gc531 (wc531, n_14068);
  nand g40927 (n_14139, n_18200, n_20856);
  nand g40928 (n_14397, n_16427, n_16428);
  or g40929 (n_18446, \data_stack_mem[4] [2], wc532);
  not gc532 (wc532, n_14022);
  or g40930 (n_19718, n_13942, wc533);
  not gc533 (wc533, n_14133);
  nand g40931 (n_21987, n_13987, n_13990);
  or g40932 (n_21988, n_13987, n_13990);
  nand g40933 (n_13991, n_21987, n_21988);
  or g40934 (n_20171, n_13942, wc534);
  not gc534 (wc534, n_14337);
  or g40935 (n_18322, \data_stack_mem[5] [1], wc535);
  not gc535 (wc535, n_13930);
  nand g40936 (n_18206, \data_stack_mem[2] [4], n_14197);
  or g40937 (n_16396, n_16395, wc536);
  not gc536 (wc536, n_13920);
  nand g40938 (n_14022, n_18194, n_20853);
  or g40939 (n_18315, wc537, n_15370);
  not gc537 (wc537, n_14032);
  or g40940 (n_18314, n_14032, wc538);
  not gc538 (wc538, n_15370);
  nand g40941 (n_16314, n_16312, n_16313);
  nand g40942 (n_14175, n_18116, n_20847);
  or g40943 (n_14055, wc539, n_18273);
  not gc539 (wc539, n_18272);
  or g40944 (n_14217, wc540, n_18258);
  not gc540 (wc540, n_18257);
  nand g40945 (n_16302, n_16300, n_16301);
  or g40946 (n_14062, wc541, n_18201);
  not gc541 (wc541, n_13914);
  nand g40947 (n_16407, n_14378, n_14425);
  or g40948 (n_16421, wc542, n_14425);
  not gc542 (wc542, n_15468);
  or g40949 (n_16408, n_14380, n_14425);
  nand g40950 (n_14068, n_18188, n_20850);
  or g40951 (n_18387, sh_reg_in[1], n_14285);
  or g40952 (n_16395, wc543, n_14379);
  not gc543 (wc543, n_14378);
  or g40953 (n_14133, wc544, n_18288);
  not gc544 (wc544, n_18287);
  nand g40954 (n_18375, n_18372, n_18373);
  or g40955 (n_16397, wc545, n_14380);
  not gc545 (wc545, n_14379);
  nand g40956 (n_18389, n_15488, sh_reg_in[1]);
  or g40957 (n_13969, n_13918, n_18189);
  or g40958 (n_18183, \data_stack_mem[3] [2], wc546);
  not gc546 (wc546, n_14032);
  or g40959 (n_18176, wc547, n_14109);
  not gc547 (wc547, n_15379);
  or g40960 (n_18177, n_15379, wc548);
  not gc548 (wc548, n_14109);
  or g40961 (n_18485, n_14246, n_14241);
  nand g40962 (n_16427, n_15469, n_14379);
  or g40963 (n_14337, wc549, n_18237);
  not gc549 (wc549, n_18236);
  nand g40964 (n_14197, n_18110, n_20844);
  nand g40965 (n_20856, n_14978, n_14066);
  nand g40966 (n_18416, n_14951, n_13929);
  or g40967 (n_14471, wc550, n_18303);
  not gc550 (wc550, n_18302);
  or g40968 (n_18170, wc551, n_14141);
  not gc551 (wc551, n_15368);
  or g40969 (n_18171, n_15368, wc552);
  not gc552 (wc552, n_14141);
  or g40970 (n_13987, n_13918, n_18195);
  nand g40971 (n_14379, n_15708, n_20823);
  nand g40972 (n_18374, n_15479, sh_reg_in[1]);
  nand g40973 (n_18195, n_14974, n_18194);
  nand g40974 (n_18189, n_15031, n_18188);
  nand g40975 (n_18258, n_18255, n_18256);
  nand g40976 (n_20844, n_14981, n_14141);
  or g40977 (n_14755, n_17276, n_17277);
  or g40978 (n_14752, n_17132, n_17133);
  nand g40979 (n_15488, n_18308, n_18309);
  or g40980 (n_14768, n_17900, n_17901);
  or g40981 (n_14760, n_17468, n_17469);
  nand g40982 (n_18288, n_18285, n_18286);
  or g40983 (n_14772, n_18092, n_18093);
  nand g40984 (n_14032, n_16439, n_16440);
  or g40985 (n_14764, n_17612, n_17613);
  or g40986 (n_14285, n_16059, wc553);
  not gc553 (wc553, n_14252);
  or g40987 (n_14770, n_17996, n_17997);
  nand g40988 (n_14066, n_16415, n_16416);
  or g40989 (n_14753, n_17180, n_17181);
  or g40990 (n_16312, n_16311, wc554);
  not gc554 (wc554, n_13920);
  nand g40991 (n_20847, n_14982, n_14109);
  nand g40992 (n_18237, n_18234, n_18235);
  nand g40993 (n_19029, n_19026, n_19027);
  or g40994 (n_14757, n_17324, n_17325);
  or g40995 (n_14767, n_17756, n_17757);
  nand g40996 (n_18303, n_18300, n_18301);
  nand g40997 (n_20853, n_14974, n_13990);
  or g40998 (n_16301, n_16299, wc555);
  not gc555 (wc555, n_13920);
  or g40999 (n_14761, n_17516, n_17517);
  nand g41000 (n_15368, n_16373, n_16374);
  nand g41001 (n_18273, n_18270, n_18271);
  nand g41002 (n_15370, n_18140, n_18141);
  or g41003 (n_14763, n_17852, n_17853);
  or g41004 (n_14246, wc556, n_16209);
  not gc556 (wc556, n_14872);
  or g41005 (n_14758, n_17372, n_17373);
  or g41006 (n_14765, n_17660, n_17661);
  or g41007 (n_18372, sh_reg_in[1], n_14009);
  nand g41008 (n_14425, n_15627, n_20820);
  or g41009 (n_14754, n_17228, n_17229);
  or g41010 (n_14769, n_17948, n_17949);
  or g41011 (n_14263, wc557, n_16185);
  not gc557 (wc557, n_14872);
  nand g41012 (n_20850, n_15031, n_13980);
  or g41013 (n_14762, n_17564, n_17565);
  or g41014 (n_14756, n_17804, n_17805);
  nand g41015 (n_15379, n_16379, n_16380);
  or g41016 (n_14759, n_17420, n_17421);
  nand g41017 (n_13929, n_18164, n_18165);
  or g41018 (n_14771, n_18044, n_18045);
  nand g41019 (n_18201, n_14978, n_18200);
  or g41020 (n_14766, n_17708, n_17709);
  or g41021 (n_18255, n_13937, n_18254);
  or g41022 (n_14703, n_17084, n_17085);
  nand g41023 (n_20823, n_15458, n_14345);
  or g41024 (n_17133, n_17130, n_17131);
  or g41025 (n_17181, n_17178, n_17179);
  or g41026 (n_18165, n_13928, n_13918);
  or g41027 (n_18308, sh_reg_in[0], wc558);
  not gc558 (wc558, n_14283);
  or g41028 (n_18116, \data_stack_mem[2] [3], wc559);
  not gc559 (wc559, n_14110);
  or g41029 (n_19026, sh_reg_in[0], wc560);
  not gc560 (wc560, n_13946);
  or g41030 (n_17229, n_17226, n_17227);
  or g41031 (n_18270, n_13937, n_18269);
  or g41032 (n_16059, n_16058, wc561);
  not gc561 (wc561, n_14234);
  nand g41033 (n_18110, \data_stack_mem[2] [3], n_14142);
  or g41034 (n_18388, n_18386, wc562);
  not gc562 (wc562, \data_stack_mem[8] [5]);
  or g41035 (n_16313, n_14311, wc563);
  not gc563 (wc563, n_14345);
  or g41036 (n_16311, wc564, n_14345);
  not gc564 (wc564, n_14310);
  or g41037 (n_18285, n_13937, n_18284);
  or g41038 (n_17277, n_17274, n_17275);
  or g41039 (n_17325, n_17322, n_17323);
  or g41040 (n_18188, wc565, n_13968);
  not gc565 (wc565, \data_stack_mem[4] [1]);
  or g41041 (n_17373, n_17370, n_17371);
  nand g41042 (n_16299, n_14310, n_14313);
  or g41043 (n_16300, n_14311, n_14313);
  or g41044 (n_17421, n_17418, n_17419);
  or g41045 (n_18300, n_13937, n_18299);
  nand g41046 (n_13980, n_18158, n_18159);
  or g41047 (n_18373, n_18371, wc566);
  not gc566 (wc566, \data_stack_mem[8] [1]);
  or g41048 (n_17469, n_17466, n_17467);
  or g41049 (n_14009, n_15978, wc567);
  not gc567 (wc567, n_13983);
  or g41050 (n_18301, sh_reg_in[0], wc568);
  not gc568 (wc568, n_14470);
  or g41051 (n_18194, \data_stack_mem[4] [1], wc569);
  not gc569 (wc569, n_13928);
  nand g41052 (n_16185, n_16183, n_16184);
  or g41053 (n_17517, n_17514, n_17515);
  or g41054 (n_17565, n_17562, n_17563);
  or g41055 (n_16374, n_14104, wc570);
  not gc570 (wc570, n_14142);
  nand g41056 (n_13990, n_18152, n_18153);
  or g41057 (n_16373, n_14103, n_14142);
  or g41058 (n_16439, wc571, n_14031);
  not gc571 (wc571, n_15342);
  or g41059 (n_17613, n_17610, n_17611);
  or g41060 (n_16440, n_15342, wc572);
  not gc572 (wc572, n_14031);
  nand g41061 (n_15479, n_18242, n_18243);
  or g41062 (n_17661, n_17658, n_17659);
  or g41063 (n_18234, n_13937, n_18233);
  or g41064 (n_17709, n_17706, n_17707);
  or g41065 (n_18140, n_14889, n_14023);
  or g41066 (n_17757, n_17754, n_17755);
  or g41067 (n_18141, n_14046, wc573);
  not gc573 (wc573, n_14023);
  or g41068 (n_18093, n_18090, n_18091);
  or g41069 (n_17805, n_17802, n_17803);
  or g41070 (n_16380, n_14103, wc574);
  not gc574 (wc574, n_14110);
  or g41071 (n_16379, n_14104, n_14110);
  or g41072 (n_17853, n_17850, n_17851);
  nand g41073 (n_20820, n_14989, n_14313);
  or g41074 (n_17901, n_17898, n_17899);
  or g41075 (n_18045, n_18042, n_18043);
  or g41076 (n_17949, n_17946, n_17947);
  nand g41077 (n_16209, n_16207, n_16208);
  or g41078 (n_17997, n_17994, n_17995);
  nand g41079 (n_18200, \data_stack_mem[3] [2], n_14061);
  or g41080 (n_16416, n_15323, wc575);
  not gc575 (wc575, n_14065);
  or g41081 (n_16415, wc576, n_14065);
  not gc576 (wc576, n_15323);
  nand g41082 (n_13867, n_16514, n_16515);
  nand g41083 (n_15323, n_16247, n_16248);
  nand g41084 (n_13866, n_16508, n_16509);
  or g41085 (n_17996, n_17992, n_17993);
  or g41086 (n_17995, wc577, n_17991);
  not gc577 (wc577, n_17990);
  or g41087 (n_18043, wc578, n_18039);
  not gc578 (wc578, n_18038);
  or g41088 (n_16208, n_16206, wc579);
  not gc579 (wc579, n_13920);
  nand g41089 (n_13865, n_16502, n_16503);
  or g41090 (n_17948, n_17944, n_17945);
  or g41091 (n_17947, wc580, n_17943);
  not gc580 (wc580, n_17942);
  or g41092 (n_18044, n_18040, n_18041);
  or g41093 (n_17900, n_17896, n_17897);
  or g41094 (n_17899, wc581, n_17895);
  not gc581 (wc581, n_17894);
  nand g41095 (n_13864, n_16496, n_16497);
  or g41096 (n_20169, wc582, n_14356);
  not gc582 (wc582, n_15373);
  nand g41097 (n_14061, n_18104, n_20841);
  nand g41098 (n_14589, n_16568, n_16569);
  or g41099 (n_17852, n_17848, n_17849);
  nand g41100 (n_14590, n_16574, n_16575);
  or g41101 (n_17851, wc583, n_17847);
  not gc583 (wc583, n_17846);
  nand g41102 (n_14591, n_16580, n_16581);
  nand g41103 (n_14110, n_16349, n_16350);
  nand g41104 (n_14592, n_16586, n_16587);
  nand g41105 (n_13863, n_16490, n_16491);
  nand g41106 (n_14593, n_16592, n_16593);
  or g41107 (n_18091, wc584, n_18087);
  not gc584 (wc584, n_18086);
  nand g41108 (n_14594, n_16598, n_16599);
  or g41109 (n_18092, n_18088, n_18089);
  nand g41110 (n_14595, n_16604, n_16605);
  or g41111 (n_17804, n_17800, n_17801);
  nand g41112 (n_14596, n_16610, n_16611);
  or g41113 (n_17803, wc585, n_17799);
  not gc585 (wc585, n_17798);
  nand g41114 (n_14599, n_16616, n_16617);
  or g41115 (n_18235, sh_reg_in[0], wc586);
  not gc586 (wc586, n_14336);
  nand g41116 (n_13862, n_16484, n_16485);
  or g41117 (n_17756, n_17752, n_17753);
  nand g41118 (n_14600, n_16622, n_16623);
  or g41119 (n_17755, wc587, n_17751);
  not gc587 (wc587, n_17750);
  nand g41120 (n_14601, n_16628, n_16629);
  nand g41121 (n_13861, n_16478, n_16479);
  nand g41122 (n_14602, n_16634, n_16635);
  or g41123 (n_17708, n_17704, n_17705);
  or g41124 (n_18242, sh_reg_in[0], wc588);
  not gc588 (wc588, n_14007);
  or g41125 (n_18233, wc589, n_14335);
  not gc589 (wc589, \data_stack_mem[8] [6]);
  nand g41126 (n_18236, n_15475, n_14335);
  or g41127 (n_17707, wc590, n_17703);
  not gc590 (wc590, n_17702);
  nand g41128 (n_14603, n_16640, n_16641);
  nand g41129 (n_14023, n_18098, n_20838);
  nand g41130 (n_14655, n_16964, n_16965);
  or g41131 (n_17660, n_17656, n_17657);
  nand g41132 (n_14605, n_16652, n_16653);
  or g41133 (n_17659, wc591, n_17655);
  not gc591 (wc591, n_17654);
  nand g41134 (n_14606, n_16658, n_16659);
  nand g41135 (n_18243, n_15478, n_14006);
  nand g41136 (n_14611, n_16664, n_16665);
  or g41137 (n_17612, n_17608, n_17609);
  or g41138 (n_20289, wc592, n_14474);
  not gc592 (wc592, n_15301);
  or g41139 (n_17611, wc593, n_17607);
  not gc593 (wc593, n_17606);
  nand g41140 (n_14612, n_16670, n_16671);
  nand g41141 (n_14142, n_16343, n_16344);
  nand g41142 (n_14613, n_16676, n_16677);
  nand g41143 (n_13860, n_16472, n_16473);
  nand g41144 (n_14614, n_16682, n_16683);
  nand g41145 (n_15342, n_16262, n_16263);
  nand g41146 (n_14615, n_16688, n_16689);
  or g41147 (n_18153, wc594, n_15351);
  not gc594 (wc594, n_13989);
  nand g41148 (n_14616, n_16694, n_16695);
  or g41149 (n_17564, n_17560, n_17561);
  nand g41150 (n_14617, n_16700, n_16701);
  or g41151 (n_17563, wc595, n_17559);
  not gc595 (wc595, n_17558);
  nand g41152 (n_14618, n_16706, n_16707);
  or g41153 (n_16183, n_16182, wc596);
  not gc596 (wc596, n_13920);
  nand g41154 (n_14621, n_16712, n_16713);
  or g41155 (n_17516, n_17512, n_17513);
  nand g41156 (n_14622, n_16718, n_16719);
  or g41157 (n_17515, wc597, n_17511);
  not gc597 (wc597, n_17510);
  or g41158 (n_18152, n_13989, wc598);
  not gc598 (wc598, n_15351);
  or g41159 (n_14470, \data_stack_mem[0] [7], n_15948);
  or g41160 (n_15978, n_15977, wc599);
  not gc599 (wc599, n_13963);
  nand g41161 (n_14623, n_16724, n_16725);
  or g41162 (n_17468, n_17464, n_17465);
  nand g41163 (n_14624, n_16730, n_16731);
  or g41164 (n_17467, wc600, n_17463);
  not gc600 (wc600, n_17462);
  nand g41165 (n_14625, n_16736, n_16737);
  or g41166 (n_18371, n_14006, n_14867);
  or g41167 (n_18299, wc601, n_14469);
  not gc601 (wc601, \data_stack_mem[8] [7]);
  nand g41168 (n_18302, n_15483, n_14469);
  or g41169 (n_18159, wc602, n_15357);
  not gc602 (wc602, n_13979);
  nand g41170 (n_14626, n_16742, n_16743);
  or g41171 (n_17420, n_17416, n_17417);
  nand g41172 (n_14627, n_16748, n_16749);
  or g41173 (n_17419, wc603, n_17415);
  not gc603 (wc603, n_17414);
  nand g41174 (n_14628, n_16754, n_16755);
  nand g41175 (n_14313, n_15624, n_20817);
  or g41176 (n_17372, n_17368, n_17369);
  or g41177 (n_17371, wc604, n_17367);
  not gc604 (wc604, n_17366);
  or g41178 (n_18158, n_13979, wc605);
  not gc605 (wc605, n_15357);
  or g41179 (n_17324, n_17320, n_17321);
  or g41180 (n_17323, wc606, n_17319);
  not gc606 (wc606, n_17318);
  nand g41181 (n_14345, n_16190, n_16191);
  or g41182 (n_17276, n_17272, n_17273);
  nand g41183 (n_18287, n_15482, n_14131);
  or g41184 (n_18284, wc607, n_14131);
  not gc607 (wc607, \data_stack_mem[8] [3]);
  or g41185 (n_17275, wc608, n_17271);
  not gc608 (wc608, n_17270);
  or g41186 (n_14199, n_16083, wc609);
  not gc609 (wc609, n_14178);
  nand g41187 (n_18272, n_15481, n_14053);
  or g41188 (n_18269, wc610, n_14053);
  not gc610 (wc610, \data_stack_mem[8] [2]);
  or g41189 (n_18386, n_14282, n_14867);
  or g41190 (n_14180, n_16071, wc611);
  not gc611 (wc611, n_14178);
  or g41191 (n_18286, sh_reg_in[0], wc612);
  not gc612 (wc612, n_14132);
  or g41192 (n_17228, n_17224, n_17225);
  or g41193 (n_17227, wc613, n_17223);
  not gc613 (wc613, n_17222);
  or g41194 (n_16058, n_16057, n_13943);
  or g41195 (n_13946, wc614, n_16029);
  not gc614 (wc614, n_13921);
  or g41196 (n_18271, sh_reg_in[0], wc615);
  not gc615 (wc615, n_14054);
  nand g41197 (n_18309, n_15487, n_14282);
  or g41198 (n_14283, \data_stack_mem[0] [5], n_15909);
  nand g41199 (n_14632, n_16856, n_16857);
  or g41200 (n_17180, n_17176, n_17177);
  or g41201 (n_17179, wc616, n_17175);
  not gc616 (wc616, n_17174);
  nand g41202 (n_14633, n_16862, n_16863);
  or g41203 (n_19716, wc617, n_14153);
  not gc617 (wc617, n_15443);
  or g41204 (n_17132, n_17128, n_17129);
  nand g41205 (n_14634, n_16868, n_16869);
  or g41206 (n_17131, wc618, n_17127);
  not gc618 (wc618, n_17126);
  nand g41207 (n_14635, n_16874, n_16875);
  or g41208 (n_17085, n_17082, n_17083);
  or g41209 (n_17084, n_17080, n_17081);
  nand g41210 (n_14636, n_16880, n_16881);
  nand g41211 (n_14692, n_17042, n_17043);
  nand g41212 (n_14691, n_17036, n_17037);
  nand g41213 (n_14637, n_16886, n_16887);
  nand g41214 (n_14690, n_17030, n_17031);
  nand g41215 (n_14689, n_17024, n_17025);
  nand g41216 (n_14638, n_16892, n_16893);
  nand g41217 (n_14688, n_17018, n_17019);
  nand g41218 (n_18257, n_15480, n_14215);
  nand g41219 (n_14639, n_16898, n_16899);
  or g41220 (n_18254, wc619, n_14215);
  not gc619 (wc619, \data_stack_mem[8] [4]);
  nand g41221 (n_14642, n_16904, n_16905);
  nand g41222 (n_18164, n_14967, n_13927);
  nand g41223 (n_14643, n_16910, n_16911);
  nand g41224 (n_14687, n_17012, n_17013);
  nand g41225 (n_14644, n_16916, n_16917);
  nand g41226 (n_14686, n_17006, n_17007);
  nand g41227 (n_14645, n_16922, n_16923);
  nand g41228 (n_14685, n_17000, n_17001);
  nand g41229 (n_14646, n_16928, n_16929);
  nand g41230 (n_14660, n_16994, n_16995);
  nand g41231 (n_14647, n_16934, n_16935);
  or g41232 (n_18256, sh_reg_in[0], wc620);
  not gc620 (wc620, n_14216);
  nand g41233 (n_14648, n_16940, n_16941);
  nand g41234 (n_14659, n_16988, n_16989);
  nand g41235 (n_14649, n_16946, n_16947);
  or g41236 (n_19941, wc621, n_14220);
  not gc621 (wc621, n_15430);
  nand g41237 (n_14658, n_16982, n_16983);
  nand g41238 (n_14657, n_16976, n_16977);
  nand g41239 (n_14653, n_16952, n_16953);
  nand g41240 (n_14656, n_16970, n_16971);
  nand g41241 (n_14654, n_16958, n_16959);
  nand g41242 (n_14604, n_16646, n_16647);
  nand g41243 (n_16971, \data_stack_mem[4] [6], n_14652);
  nand g41244 (n_16965, \data_stack_mem[4] [7], n_14652);
  nand g41245 (n_16977, \data_stack_mem[4] [5], n_14652);
  nand g41246 (n_16959, \data_stack_mem[4] [0], n_14652);
  nand g41247 (n_16983, \data_stack_mem[4] [4], n_14652);
  nand g41248 (n_16953, \data_stack_mem[4] [2], n_14652);
  nand g41249 (n_16989, \data_stack_mem[4] [3], n_14652);
  or g41250 (n_14220, n_16047, wc622);
  not gc622 (wc622, n_14174);
  nand g41251 (n_16995, \data_stack_mem[4] [1], n_14652);
  nand g41252 (n_16947, \data_stack_mem[0] [3], n_14640);
  or g41253 (n_14216, \data_stack_mem[0] [4], n_15888);
  nand g41254 (n_16941, \data_stack_mem[0] [2], n_14640);
  nand g41255 (n_17001, \data_stack_mem[5] [7], n_14684);
  nand g41256 (n_16935, \data_stack_mem[0] [1], n_14640);
  nand g41257 (n_17007, \data_stack_mem[5] [6], n_14684);
  nand g41258 (n_16929, \data_stack_mem[0] [0], n_14640);
  nand g41259 (n_17013, \data_stack_mem[5] [5], n_14684);
  nand g41260 (n_16923, \data_stack_mem[0] [5], n_14640);
  nand g41261 (n_16917, \data_stack_mem[0] [7], n_14640);
  nand g41262 (n_16911, \data_stack_mem[0] [4], n_14640);
  nand g41263 (n_16905, \data_stack_mem[0] [6], n_14640);
  nand g41264 (n_17019, \data_stack_mem[5] [4], n_14684);
  nand g41265 (n_16899, \data_stack_mem[1] [0], n_14630);
  nand g41266 (n_17025, \data_stack_mem[5] [3], n_14684);
  or g41267 (n_16898, wc623, n_14631);
  not gc623 (wc623, sh_reg_in[0]);
  nand g41268 (n_17031, \data_stack_mem[5] [1], n_14684);
  nand g41269 (n_16893, \data_stack_mem[1] [1], n_14630);
  nand g41270 (n_17037, \data_stack_mem[5] [2], n_14684);
  or g41271 (n_16892, wc624, n_14631);
  not gc624 (wc624, sh_reg_in[1]);
  nand g41272 (n_17043, \data_stack_mem[5] [0], n_14684);
  nand g41273 (n_16887, \data_stack_mem[1] [2], n_14630);
  nand g41274 (n_17080, n_17072, n_17073);
  nand g41275 (n_17081, n_17074, n_17075);
  nand g41276 (n_17082, n_17076, n_17077);
  nand g41277 (n_17083, n_17078, n_17079);
  or g41278 (n_16886, wc625, n_14631);
  not gc625 (wc625, sh_reg_in[2]);
  nand g41279 (n_16881, \data_stack_mem[1] [3], n_14630);
  or g41280 (n_16880, wc626, n_14631);
  not gc626 (wc626, sh_reg_in[3]);
  nand g41281 (n_17127, n_17118, n_17119);
  nand g41282 (n_17128, n_17120, n_17121);
  nand g41283 (n_17129, n_17122, n_17123);
  or g41284 (n_19563, wc627, n_14076);
  not gc627 (wc627, n_15447);
  nand g41285 (n_17130, n_17124, n_17125);
  nand g41286 (n_16875, \data_stack_mem[1] [4], n_14630);
  or g41287 (n_16874, wc628, n_14631);
  not gc628 (wc628, sh_reg_in[4]);
  nand g41288 (n_16869, \data_stack_mem[1] [5], n_14630);
  nand g41289 (n_17175, n_17166, n_17167);
  nand g41290 (n_17176, n_17168, n_17169);
  nand g41291 (n_17177, n_17170, n_17171);
  nand g41292 (n_17178, n_17172, n_17173);
  or g41293 (n_16868, wc629, n_14631);
  not gc629 (wc629, sh_reg_in[5]);
  nand g41294 (n_16863, \data_stack_mem[1] [6], n_14630);
  or g41295 (n_16862, wc630, n_14631);
  not gc630 (wc630, sh_reg_in[6]);
  nand g41296 (n_16857, \data_stack_mem[1] [7], n_14630);
  or g41297 (n_16856, wc631, n_14631);
  not gc631 (wc631, sh_reg_in[7]);
  nand g41298 (n_17223, n_17214, n_17215);
  nand g41299 (n_17224, n_17216, n_17217);
  nand g41300 (n_17225, n_17218, n_17219);
  nand g41301 (n_14576, n_16850, n_16851);
  or g41302 (n_14054, \data_stack_mem[0] [2], n_15846);
  nand g41303 (n_17226, n_17220, n_17221);
  or g41304 (n_16029, n_16028, wc632);
  not gc632 (wc632, n_14980);
  nand g41305 (n_14574, n_16844, n_16845);
  nand g41306 (n_14572, n_16838, n_16839);
  nand g41307 (n_14570, n_16832, n_16833);
  nand g41308 (n_16071, n_16069, n_16070);
  nand g41309 (n_14568, n_16826, n_16827);
  nand g41310 (n_14566, n_16820, n_16821);
  nand g41311 (n_14564, n_16814, n_16815);
  nand g41312 (n_17271, n_17262, n_17263);
  nand g41313 (n_17272, n_17264, n_17265);
  nand g41314 (n_17273, n_17266, n_17267);
  nand g41315 (n_17274, n_17268, n_17269);
  nand g41316 (n_16083, n_16081, n_16082);
  nand g41317 (n_14562, n_16808, n_16809);
  nand g41318 (n_13901, n_16802, n_16803);
  nand g41319 (n_17319, n_17310, n_17311);
  nand g41320 (n_17320, n_17312, n_17313);
  nand g41321 (n_17321, n_17314, n_17315);
  nand g41322 (n_17322, n_17316, n_17317);
  nand g41323 (n_13898, n_16796, n_16797);
  nand g41324 (n_13895, n_16790, n_16791);
  nand g41325 (n_13892, n_16784, n_16785);
  nand g41326 (n_17367, n_17358, n_17359);
  nand g41327 (n_17368, n_17360, n_17361);
  nand g41328 (n_17369, n_17362, n_17363);
  nand g41329 (n_17370, n_17364, n_17365);
  nand g41330 (n_13889, n_16778, n_16779);
  nand g41331 (n_13886, n_16772, n_16773);
  nand g41332 (n_13883, n_16766, n_16767);
  nand g41333 (n_17415, n_17406, n_17407);
  nand g41334 (n_17416, n_17408, n_17409);
  nand g41335 (n_17417, n_17410, n_17411);
  nand g41336 (n_17418, n_17412, n_17413);
  nand g41337 (n_13880, n_16760, n_16761);
  nand g41338 (n_16755, \data_stack_mem[6] [7], n_14620);
  nand g41339 (n_16749, \data_stack_mem[6] [6], n_14620);
  nand g41340 (n_17463, n_17454, n_17455);
  nand g41341 (n_17464, n_17456, n_17457);
  nand g41342 (n_17465, n_17458, n_17459);
  nand g41343 (n_17466, n_17460, n_17461);
  nand g41344 (n_16743, \data_stack_mem[6] [5], n_14620);
  nand g41345 (n_16737, \data_stack_mem[6] [4], n_14620);
  nand g41346 (n_16731, \data_stack_mem[6] [3], n_14620);
  nand g41347 (n_17511, n_17502, n_17503);
  nand g41348 (n_17512, n_17504, n_17505);
  nand g41349 (n_17513, n_17506, n_17507);
  nand g41350 (n_17514, n_17508, n_17509);
  or g41351 (n_15948, wc633, n_15947);
  not gc633 (wc633, n_14396);
  nand g41352 (n_16725, \data_stack_mem[6] [2], n_14620);
  nand g41353 (n_16719, \data_stack_mem[6] [1], n_14620);
  nand g41354 (n_17559, n_17550, n_17551);
  nand g41355 (n_17560, n_17552, n_17553);
  nand g41356 (n_17561, n_17554, n_17555);
  nand g41357 (n_17562, n_17556, n_17557);
  nand g41358 (n_16713, \data_stack_mem[6] [0], n_14620);
  nand g41359 (n_16707, \data_stack_mem[7] [6], n_14610);
  nand g41360 (n_16701, \data_stack_mem[7] [3], n_14610);
  nand g41361 (n_16695, \data_stack_mem[7] [4], n_14610);
  nand g41362 (n_16689, \data_stack_mem[7] [2], n_14610);
  nand g41363 (n_16683, \data_stack_mem[7] [1], n_14610);
  nand g41364 (n_16343, n_15330, n_14063);
  nand g41365 (n_17607, n_17598, n_17599);
  nand g41366 (n_17608, n_17600, n_17601);
  nand g41367 (n_17609, n_17602, n_17603);
  nand g41368 (n_17610, n_17604, n_17605);
  nand g41369 (n_16677, \data_stack_mem[7] [7], n_14610);
  or g41370 (n_14474, n_16155, wc634);
  not gc634 (wc634, n_14411);
  nand g41371 (n_16671, \data_stack_mem[7] [0], n_14610);
  nand g41372 (n_17655, n_17646, n_17647);
  nand g41373 (n_17656, n_17648, n_17649);
  nand g41374 (n_17657, n_17650, n_17651);
  nand g41375 (n_17658, n_17652, n_17653);
  nand g41376 (n_16665, \data_stack_mem[7] [5], n_14610);
  nand g41377 (n_16659, \data_stack_mem[3] [5], n_14598);
  nand g41378 (n_16653, \data_stack_mem[3] [2], n_14598);
  nand g41379 (n_21989, n_14094, n_14130);
  or g41380 (n_21990, n_14094, n_14130);
  nand g41381 (n_14131, n_21989, n_21990);
  nand g41382 (n_17703, n_17694, n_17695);
  nand g41383 (n_17704, n_17696, n_17697);
  nand g41384 (n_17705, n_17698, n_17699);
  nand g41385 (n_17706, n_17700, n_17701);
  nand g41386 (n_16647, \data_stack_mem[3] [1], n_14598);
  nand g41387 (n_16641, \data_stack_mem[3] [7], n_14598);
  nand g41388 (n_21991, n_14208, n_14214);
  or g41389 (n_21992, n_14208, n_14214);
  nand g41390 (n_14215, n_21991, n_21992);
  nand g41391 (n_17751, n_17742, n_17743);
  nand g41392 (n_17752, n_17744, n_17745);
  nand g41393 (n_17753, n_17746, n_17747);
  nand g41394 (n_17754, n_17748, n_17749);
  nand g41395 (n_16635, \data_stack_mem[3] [4], n_14598);
  nand g41396 (n_16629, \data_stack_mem[3] [3], n_14598);
  nand g41397 (n_16623, \data_stack_mem[3] [0], n_14598);
  nand g41398 (n_17799, n_17790, n_17791);
  nand g41399 (n_17800, n_17792, n_17793);
  nand g41400 (n_17801, n_17794, n_17795);
  nand g41401 (n_17802, n_17796, n_17797);
  or g41402 (n_14336, \data_stack_mem[0] [6], n_15930);
  nand g41403 (n_16617, \data_stack_mem[3] [6], n_14598);
  nand g41404 (n_16611, \data_stack_mem[2] [7], n_14588);
  nand g41405 (n_16605, \data_stack_mem[2] [0], n_14588);
  nand g41406 (n_16599, \data_stack_mem[2] [1], n_14588);
  nand g41407 (n_16593, \data_stack_mem[2] [2], n_14588);
  nand g41408 (n_16349, n_15377, n_14026);
  nand g41409 (n_17847, n_17838, n_17839);
  nand g41410 (n_21993, n_14410, n_14468);
  or g41411 (n_21994, n_14410, n_14468);
  nand g41412 (n_14469, n_21993, n_21994);
  nand g41413 (n_17848, n_17840, n_17841);
  nand g41414 (n_17849, n_17842, n_17843);
  nand g41415 (n_17850, n_17844, n_17845);
  nand g41416 (n_16587, \data_stack_mem[2] [3], n_14588);
  nand g41417 (n_16581, \data_stack_mem[2] [6], n_14588);
  nand g41418 (n_16575, \data_stack_mem[2] [5], n_14588);
  or g41419 (n_14356, n_16152, wc635);
  not gc635 (wc635, n_14322);
  nand g41420 (n_17895, n_17886, n_17887);
  nand g41421 (n_17896, n_17888, n_17889);
  nand g41422 (n_17897, n_17890, n_17891);
  nand g41423 (n_17898, n_17892, n_17893);
  nand g41424 (n_16569, \data_stack_mem[2] [4], n_14588);
  nand g41425 (n_14577, n_16562, n_16563);
  nand g41426 (n_14575, n_16556, n_16557);
  nand g41427 (n_17943, n_17934, n_17935);
  nand g41428 (n_17944, n_17936, n_17937);
  nand g41429 (n_17945, n_17938, n_17939);
  nand g41430 (n_17946, n_17940, n_17941);
  nand g41431 (n_14573, n_16550, n_16551);
  or g41432 (n_16207, n_14244, n_14245);
  nand g41433 (n_16206, n_14243, n_14245);
  nand g41434 (n_17991, n_17982, n_17983);
  nand g41435 (n_17992, n_17984, n_17985);
  nand g41436 (n_17993, n_17986, n_17987);
  nand g41437 (n_17994, n_17988, n_17989);
  nand g41438 (n_14571, n_16544, n_16545);
  nand g41439 (n_14569, n_16538, n_16539);
  nand g41440 (n_14567, n_16532, n_16533);
  nand g41441 (n_14565, n_16526, n_16527);
  nand g41442 (n_14563, n_16520, n_16521);
  nand g41443 (n_16515, \data_stack_mem[8] [4], n_13857);
  or g41444 (n_16248, n_14025, wc636);
  not gc636 (wc636, n_14063);
  or g41445 (n_16247, n_14024, n_14063);
  or g41446 (n_16514, wc637, n_13859);
  not gc637 (wc637, sh_reg_in[4]);
  nand g41447 (n_18039, n_18030, n_18031);
  nand g41448 (n_18040, n_18032, n_18033);
  nand g41449 (n_18041, n_18034, n_18035);
  nand g41450 (n_18042, n_18036, n_18037);
  nand g41451 (n_16509, \data_stack_mem[8] [0], n_13857);
  or g41452 (n_16508, wc638, n_13859);
  not gc638 (wc638, sh_reg_in[0]);
  nand g41453 (n_16503, \data_stack_mem[8] [2], n_13857);
  or g41454 (n_16502, wc639, n_13859);
  not gc639 (wc639, sh_reg_in[2]);
  nand g41455 (n_16497, \data_stack_mem[8] [1], n_13857);
  nand g41456 (n_20841, n_14983, n_13979);
  nand g41457 (n_18087, n_18078, n_18079);
  nand g41458 (n_18088, n_18080, n_18081);
  nand g41459 (n_18089, n_18082, n_18083);
  nand g41460 (n_18090, n_18084, n_18085);
  or g41461 (n_16496, wc640, n_13859);
  not gc640 (wc640, sh_reg_in[1]);
  nand g41462 (n_16491, \data_stack_mem[8] [3], n_13857);
  or g41463 (n_16490, wc641, n_13859);
  not gc641 (wc641, sh_reg_in[3]);
  nand g41464 (n_21995, n_14015, n_14052);
  or g41465 (n_21996, n_14015, n_14052);
  nand g41466 (n_14053, n_21995, n_21996);
  nand g41467 (n_16485, \data_stack_mem[8] [6], n_13857);
  or g41468 (n_16484, wc642, n_13859);
  not gc642 (wc642, sh_reg_in[6]);
  or g41469 (n_14007, \data_stack_mem[0] [1], n_15825);
  nand g41470 (n_20838, n_14930, n_13989);
  nand g41471 (n_16479, \data_stack_mem[8] [5], n_13857);
  or g41472 (n_16478, wc643, n_13859);
  not gc643 (wc643, sh_reg_in[5]);
  nand g41473 (n_16473, \data_stack_mem[8] [7], n_13857);
  or g41474 (n_16263, n_14024, wc644);
  not gc644 (wc644, n_14026);
  or g41475 (n_16262, n_14025, n_14026);
  nand g41476 (n_21997, n_13962, n_14005);
  or g41477 (n_21998, n_13962, n_14005);
  nand g41478 (n_14006, n_21997, n_21998);
  or g41479 (n_16472, wc645, n_13859);
  not gc645 (wc645, sh_reg_in[7]);
  nand g41480 (n_14681, n_16280, n_14609);
  or g41481 (n_16182, wc646, n_14262);
  not gc646 (wc646, n_14243);
  nand g41482 (n_15351, n_16361, n_16362);
  or g41483 (n_16184, n_14244, wc647);
  not gc647 (wc647, n_14262);
  or g41484 (n_15977, n_15976, n_13943);
  nand g41485 (n_21999, n_14233, n_14281);
  or g41486 (n_22000, n_14233, n_14281);
  nand g41487 (n_14282, n_21999, n_22000);
  nand g41490 (n_20817, n_14995, n_14245);
  nand g41491 (n_15357, n_16367, n_16368);
  nand g41492 (n_22002, n_14298, n_14334);
  or g41493 (n_22003, n_14298, n_14334);
  nand g41494 (n_14335, n_22002, n_22003);
  nand g41495 (n_16190, n_15451, n_14262);
  or g41496 (n_14132, \data_stack_mem[0] [3], n_15867);
  or g41497 (n_16057, n_16056, wc648);
  not gc648 (wc648, n_14877);
  or g41498 (n_15909, n_15908, wc649);
  not gc649 (wc649, n_14240);
  or g41499 (n_14153, n_16158, wc650);
  not gc650 (wc650, n_14118);
  nand g41500 (n_13927, n_16433, n_16434);
  or g41501 (n_16610, wc651, n_14584);
  not gc651 (wc651, sh_reg_in[7]);
  or g41502 (n_16616, wc652, n_14597);
  not gc652 (wc652, sh_reg_in[6]);
  or g41503 (n_16622, wc653, n_14597);
  not gc653 (wc653, sh_reg_in[0]);
  or g41504 (n_16628, wc654, n_14597);
  not gc654 (wc654, sh_reg_in[3]);
  or g41505 (n_19260, wc655, n_13887);
  not gc655 (wc655, \out_fifo[6][0] [1]);
  or g41506 (n_19266, wc656, n_13890);
  not gc656 (wc656, \out_fifo[3][0] [1]);
  or g41507 (n_19272, wc657, n_13893);
  not gc657 (wc657, \out_fifo[7][0] [1]);
  or g41508 (n_16634, wc658, n_14597);
  not gc658 (wc658, sh_reg_in[4]);
  nand g41509 (n_22004, n_14166, n_14213);
  or g41510 (n_22005, n_14166, n_14213);
  nand g41511 (n_14214, n_22004, n_22005);
  or g41512 (n_19278, wc659, n_13896);
  not gc659 (wc659, \out_fifo[0][0] [1]);
  or g41513 (n_19284, wc660, n_13899);
  not gc660 (wc660, \out_fifo[4][0] [1]);
  nand g41514 (n_22006, n_14044, n_14051);
  or g41515 (n_22007, n_14044, n_14051);
  nand g41516 (n_14052, n_22006, n_22007);
  nand g41517 (n_22008, n_14461, n_14467);
  or g41518 (n_22009, n_14461, n_14467);
  nand g41519 (n_14468, n_22008, n_22009);
  or g41520 (n_20361, wc661, n_13881);
  not gc661 (wc661, \out_fifo[2][0] [8]);
  or g41521 (n_20466, wc662, n_13899);
  not gc662 (wc662, \out_fifo[4][1] [8]);
  or g41522 (n_20463, wc663, n_13899);
  not gc663 (wc663, \out_fifo[4][1] [6]);
  or g41523 (n_20226, wc664, n_13887);
  not gc664 (wc664, \out_fifo[6][0] [7]);
  or g41524 (n_16640, wc665, n_14597);
  not gc665 (wc665, sh_reg_in[7]);
  or g41525 (n_16646, wc666, n_14597);
  not gc666 (wc666, sh_reg_in[1]);
  or g41526 (n_16652, wc667, n_14597);
  not gc667 (wc667, sh_reg_in[2]);
  or g41527 (n_16658, wc668, n_14597);
  not gc668 (wc668, sh_reg_in[5]);
  or g41528 (n_16664, wc669, n_14609);
  not gc669 (wc669, sh_reg_in[5]);
  or g41529 (n_16670, wc670, n_14609);
  not gc670 (wc670, sh_reg_in[0]);
  or g41530 (n_15846, n_15845, wc671);
  not gc671 (wc671, n_14024);
  or g41531 (n_16676, wc672, n_14609);
  not gc672 (wc672, sh_reg_in[7]);
  or g41532 (n_16682, wc673, n_14609);
  not gc673 (wc673, sh_reg_in[1]);
  or g41533 (n_16688, wc674, n_14609);
  not gc674 (wc674, sh_reg_in[2]);
  or g41534 (n_16694, wc675, n_14609);
  not gc675 (wc675, sh_reg_in[4]);
  or g41535 (n_16700, wc676, n_14609);
  not gc676 (wc676, sh_reg_in[3]);
  or g41536 (n_16706, wc677, n_14609);
  not gc677 (wc677, sh_reg_in[6]);
  or g41537 (n_16712, wc678, n_14619);
  not gc678 (wc678, sh_reg_in[0]);
  or g41538 (n_16718, wc679, n_14619);
  not gc679 (wc679, sh_reg_in[1]);
  or g41539 (n_16724, wc680, n_14619);
  not gc680 (wc680, sh_reg_in[2]);
  or g41540 (n_16730, wc681, n_14619);
  not gc681 (wc681, sh_reg_in[3]);
  or g41541 (n_16736, wc682, n_14619);
  not gc682 (wc682, sh_reg_in[4]);
  or g41542 (n_16742, wc683, n_14619);
  not gc683 (wc683, sh_reg_in[5]);
  or g41543 (n_16748, wc684, n_14619);
  not gc684 (wc684, sh_reg_in[6]);
  or g41544 (n_16754, wc685, n_14619);
  not gc685 (wc685, sh_reg_in[7]);
  or g41545 (n_14076, n_16167, wc686);
  not gc686 (wc686, n_14037);
  or g41546 (n_16760, n_13877, n_13879);
  or g41547 (n_16761, wc687, n_13878);
  not gc687 (wc687, \out_fifo[5][2] [0]);
  or g41548 (n_16766, n_13877, n_13882);
  or g41549 (n_16767, wc688, n_13881);
  not gc688 (wc688, \out_fifo[2][2] [0]);
  or g41550 (n_16772, n_13877, n_13885);
  or g41551 (n_16773, wc689, n_13884);
  not gc689 (wc689, \out_fifo[1][2] [0]);
  or g41552 (n_16778, n_13877, n_13888);
  or g41553 (n_16779, wc690, n_13887);
  not gc690 (wc690, \out_fifo[6][2] [0]);
  or g41554 (n_16784, n_13877, n_13891);
  or g41555 (n_16785, wc691, n_13890);
  not gc691 (wc691, \out_fifo[3][2] [0]);
  or g41556 (n_16790, n_13877, n_13894);
  or g41557 (n_16791, wc692, n_13893);
  not gc692 (wc692, \out_fifo[7][2] [0]);
  or g41558 (n_16796, n_13877, n_13897);
  or g41559 (n_16797, wc693, n_13896);
  not gc693 (wc693, \out_fifo[0][2] [0]);
  or g41560 (n_15888, n_15887, wc694);
  not gc694 (wc694, n_14173);
  or g41561 (n_16802, n_13877, n_13900);
  or g41562 (n_16803, wc695, n_13899);
  not gc695 (wc695, \out_fifo[4][2] [0]);
  or g41563 (n_16808, n_13870, n_13879);
  or g41564 (n_16809, wc696, n_13878);
  not gc696 (wc696, \out_fifo[5][2] [1]);
  or g41565 (n_16814, n_13870, n_13882);
  or g41566 (n_16082, n_16080, wc697);
  not gc697 (wc697, n_13920);
  or g41567 (n_20502, wc698, n_13884);
  not gc698 (wc698, \out_fifo[1][1] [6]);
  or g41568 (n_20232, wc699, n_13890);
  not gc699 (wc699, \out_fifo[3][0] [7]);
  or g41569 (n_20499, wc700, n_13884);
  not gc700 (wc700, \out_fifo[1][1] [8]);
  or g41570 (n_16047, n_16046, wc701);
  not gc701 (wc701, n_14171);
  or g41571 (n_20238, wc702, n_13893);
  not gc702 (wc702, \out_fifo[7][0] [7]);
  or g41572 (n_20496, wc703, n_13884);
  not gc703 (wc703, \out_fifo[1][1] [7]);
  or g41573 (n_20244, wc704, n_13896);
  not gc704 (wc704, \out_fifo[0][0] [7]);
  or g41574 (n_16815, wc705, n_13881);
  not gc705 (wc705, \out_fifo[2][2] [1]);
  or g41575 (n_16820, n_13870, n_13885);
  or g41576 (n_16821, wc706, n_13884);
  not gc706 (wc706, \out_fifo[1][2] [1]);
  or g41577 (n_16826, n_13870, n_13888);
  or g41578 (n_16827, wc707, n_13887);
  not gc707 (wc707, \out_fifo[6][2] [1]);
  or g41579 (n_16832, n_13870, n_13891);
  or g41580 (n_16833, wc708, n_13890);
  not gc708 (wc708, \out_fifo[3][2] [1]);
  or g41581 (n_16838, n_13870, n_13894);
  or g41582 (n_16839, wc709, n_13893);
  not gc709 (wc709, \out_fifo[7][2] [1]);
  or g41583 (n_16844, n_13870, n_13897);
  or g41584 (n_16845, wc710, n_13896);
  not gc710 (wc710, \out_fifo[0][2] [1]);
  or g41585 (n_16850, n_13870, n_13900);
  or g41586 (n_16851, wc711, n_13899);
  not gc711 (wc711, \out_fifo[4][2] [1]);
  or g41587 (n_20493, wc712, n_13893);
  not gc712 (wc712, \out_fifo[7][1] [6]);
  or g41588 (n_19153, wc713, n_13950);
  not gc713 (wc713, n_15455);
  or g41589 (n_14631, n_20832, wc714);
  not gc714 (wc714, data_stack_pointer[0]);
  or g41590 (n_16904, wc715, n_14641);
  not gc715 (wc715, sh_reg_in[6]);
  or g41591 (n_16910, wc716, n_14641);
  not gc716 (wc716, sh_reg_in[4]);
  or g41592 (n_16916, wc717, n_14641);
  not gc717 (wc717, sh_reg_in[7]);
  or g41593 (n_16922, wc718, n_14641);
  not gc718 (wc718, sh_reg_in[5]);
  or g41594 (n_16928, wc719, n_14641);
  not gc719 (wc719, sh_reg_in[0]);
  or g41595 (n_16028, n_16027, wc720);
  not gc720 (wc720, n_15022);
  or g41596 (n_16934, wc721, n_14641);
  not gc721 (wc721, sh_reg_in[1]);
  or g41597 (n_16940, wc722, n_14641);
  not gc722 (wc722, sh_reg_in[2]);
  or g41598 (n_16946, wc723, n_14641);
  not gc723 (wc723, sh_reg_in[3]);
  or g41599 (n_20799, wc724, n_13899);
  not gc724 (wc724, \out_fifo[4][1] [0]);
  or g41600 (n_16952, wc725, n_14650);
  not gc725 (wc725, sh_reg_in[2]);
  or g41601 (n_20793, wc726, n_13896);
  not gc726 (wc726, \out_fifo[0][1] [0]);
  or g41602 (n_20787, wc727, n_13893);
  not gc727 (wc727, \out_fifo[7][1] [0]);
  or g41603 (n_19431, wc728, n_13878);
  not gc728 (wc728, \out_fifo[5][0] [2]);
  or g41604 (n_20781, wc729, n_13890);
  not gc729 (wc729, \out_fifo[3][1] [0]);
  or g41605 (n_20775, wc730, n_13887);
  not gc730 (wc730, \out_fifo[6][1] [0]);
  or g41606 (n_20769, wc731, n_13884);
  not gc731 (wc731, \out_fifo[1][1] [0]);
  nand g41607 (n_14652, n_16451, n_20835);
  or g41608 (n_16958, wc732, n_14650);
  not gc732 (wc732, sh_reg_in[0]);
  or g41609 (n_16964, wc733, n_14650);
  not gc733 (wc733, sh_reg_in[7]);
  or g41610 (n_16970, wc734, n_14650);
  not gc734 (wc734, sh_reg_in[6]);
  or g41611 (n_16976, wc735, n_14650);
  not gc735 (wc735, sh_reg_in[5]);
  or g41612 (n_16982, wc736, n_14650);
  not gc736 (wc736, sh_reg_in[4]);
  or g41613 (n_16988, wc737, n_14650);
  not gc737 (wc737, sh_reg_in[3]);
  or g41614 (n_16994, wc738, n_14650);
  not gc738 (wc738, sh_reg_in[1]);
  or g41615 (n_17000, wc739, n_14683);
  not gc739 (wc739, sh_reg_in[7]);
  or g41616 (n_17006, wc740, n_14683);
  not gc740 (wc740, sh_reg_in[6]);
  or g41617 (n_15947, n_15946, wc741);
  not gc741 (wc741, n_14410);
  or g41618 (n_17012, wc742, n_14683);
  not gc742 (wc742, sh_reg_in[5]);
  or g41619 (n_17018, wc743, n_14683);
  not gc743 (wc743, sh_reg_in[4]);
  or g41620 (n_17024, wc744, n_14683);
  not gc744 (wc744, sh_reg_in[3]);
  or g41621 (n_17030, wc745, n_14683);
  not gc745 (wc745, sh_reg_in[1]);
  or g41622 (n_17036, wc746, n_14683);
  not gc746 (wc746, sh_reg_in[2]);
  or g41623 (n_19437, wc747, n_13881);
  not gc747 (wc747, \out_fifo[2][0] [2]);
  or g41624 (n_17042, wc748, n_14683);
  not gc748 (wc748, sh_reg_in[0]);
  or g41625 (n_17072, wc749, n_14702);
  not gc749 (wc749, \out_fifo[7][0] [0]);
  or g41626 (n_19443, wc750, n_13884);
  not gc750 (wc750, \out_fifo[1][0] [2]);
  or g41627 (n_17073, wc751, n_14701);
  not gc751 (wc751, \out_fifo[3][0] [0]);
  or g41628 (n_16155, wc752, n_14473);
  not gc752 (wc752, n_15496);
  or g41629 (n_17074, wc753, n_14700);
  not gc753 (wc753, \out_fifo[5][0] [0]);
  or g41630 (n_20763, wc754, n_13881);
  not gc754 (wc754, \out_fifo[2][1] [0]);
  or g41631 (n_20757, wc755, n_13878);
  not gc755 (wc755, \out_fifo[5][1] [0]);
  or g41632 (n_20751, wc756, n_13899);
  not gc756 (wc756, \out_fifo[4][0] [0]);
  or g41633 (n_20745, wc757, n_13896);
  not gc757 (wc757, \out_fifo[0][0] [0]);
  or g41634 (n_20739, wc758, n_13893);
  not gc758 (wc758, \out_fifo[7][0] [0]);
  or g41635 (n_17075, wc759, n_14699);
  not gc759 (wc759, \out_fifo[1][0] [0]);
  or g41636 (n_17076, wc760, n_14697);
  not gc760 (wc760, \out_fifo[0][0] [0]);
  or g41637 (n_17077, wc761, n_14696);
  not gc761 (wc761, \out_fifo[2][0] [0]);
  or g41638 (n_17078, wc762, n_14695);
  not gc762 (wc762, \out_fifo[4][0] [0]);
  or g41639 (n_17079, wc763, n_14694);
  not gc763 (wc763, \out_fifo[6][0] [0]);
  or g41640 (n_17118, wc764, n_14701);
  not gc764 (wc764, \out_fifo[3][0] [8]);
  or g41641 (n_17119, wc765, n_14702);
  not gc765 (wc765, \out_fifo[7][0] [8]);
  or g41642 (n_19449, wc766, n_13887);
  not gc766 (wc766, \out_fifo[6][0] [2]);
  or g41643 (n_17120, wc767, n_14700);
  not gc767 (wc767, \out_fifo[5][0] [8]);
  or g41644 (n_15930, n_15929, wc768);
  not gc768 (wc768, n_14307);
  or g41645 (n_17121, wc769, n_14699);
  not gc769 (wc769, \out_fifo[1][0] [8]);
  or g41646 (n_19455, wc770, n_13890);
  not gc770 (wc770, \out_fifo[3][0] [2]);
  or g41647 (n_17123, wc771, n_14694);
  not gc771 (wc771, \out_fifo[6][0] [8]);
  or g41648 (n_17124, wc772, n_14695);
  not gc772 (wc772, \out_fifo[4][0] [8]);
  or g41649 (n_19461, wc773, n_13893);
  not gc773 (wc773, \out_fifo[7][0] [2]);
  or g41650 (n_17125, wc774, n_14696);
  not gc774 (wc774, \out_fifo[2][0] [8]);
  or g41651 (n_17126, wc775, n_14697);
  not gc775 (wc775, \out_fifo[0][0] [8]);
  or g41652 (n_17166, wc776, n_14701);
  not gc776 (wc776, \out_fifo[3][1] [6]);
  or g41653 (n_17167, wc777, n_14702);
  not gc777 (wc777, \out_fifo[7][1] [6]);
  or g41654 (n_17168, wc778, n_14700);
  not gc778 (wc778, \out_fifo[5][1] [6]);
  or g41655 (n_19467, wc779, n_13896);
  not gc779 (wc779, \out_fifo[0][0] [2]);
  or g41656 (n_17169, wc780, n_14699);
  not gc780 (wc780, \out_fifo[1][1] [6]);
  or g41657 (n_20367, wc781, n_13884);
  not gc781 (wc781, \out_fifo[1][1] [1]);
  or g41658 (n_16152, wc782, n_14355);
  not gc782 (wc782, n_15493);
  or g41659 (n_17171, wc783, n_14694);
  not gc783 (wc783, \out_fifo[6][1] [6]);
  or g41660 (n_17172, wc784, n_14695);
  not gc784 (wc784, \out_fifo[4][1] [6]);
  or g41661 (n_19473, wc785, n_13899);
  not gc785 (wc785, \out_fifo[4][0] [2]);
  or g41662 (n_17173, wc786, n_14696);
  not gc786 (wc786, \out_fifo[2][1] [6]);
  or g41663 (n_17174, wc787, n_14697);
  not gc787 (wc787, \out_fifo[0][1] [6]);
  or g41664 (n_17214, wc788, n_14701);
  not gc788 (wc788, \out_fifo[3][0] [7]);
  or g41665 (n_17215, wc789, n_14702);
  not gc789 (wc789, \out_fifo[7][0] [7]);
  or g41666 (n_17216, wc790, n_14700);
  not gc790 (wc790, \out_fifo[5][0] [7]);
  or g41667 (n_19644, wc791, n_13878);
  not gc791 (wc791, \out_fifo[5][0] [3]);
  or g41668 (n_17217, wc792, n_14699);
  not gc792 (wc792, \out_fifo[1][0] [7]);
  or g41669 (n_15825, n_15824, wc793);
  not gc793 (wc793, n_13973);
  or g41670 (n_19650, wc794, n_13881);
  not gc794 (wc794, \out_fifo[2][0] [3]);
  or g41671 (n_17219, wc795, n_14694);
  not gc795 (wc795, \out_fifo[6][0] [7]);
  or g41672 (n_17220, wc796, n_14695);
  not gc796 (wc796, \out_fifo[4][0] [7]);
  or g41673 (n_17221, wc797, n_14696);
  not gc797 (wc797, \out_fifo[2][0] [7]);
  or g41674 (n_20250, wc798, n_13899);
  not gc798 (wc798, \out_fifo[4][0] [7]);
  or g41675 (n_17222, wc799, n_14697);
  not gc799 (wc799, \out_fifo[0][0] [7]);
  or g41676 (n_19656, wc800, n_13884);
  not gc800 (wc800, \out_fifo[1][0] [3]);
  or g41677 (n_17262, wc801, n_14701);
  not gc801 (wc801, \out_fifo[3][1] [7]);
  or g41678 (n_19662, wc802, n_13887);
  not gc802 (wc802, \out_fifo[6][0] [3]);
  or g41679 (n_19668, wc803, n_13890);
  not gc803 (wc803, \out_fifo[3][0] [3]);
  or g41680 (n_16069, n_16068, wc804);
  not gc804 (wc804, n_13920);
  or g41681 (n_19674, wc805, n_13893);
  not gc805 (wc805, \out_fifo[7][0] [3]);
  or g41682 (n_15976, n_14008, n_15975);
  or g41683 (n_19680, wc806, n_13896);
  not gc806 (wc806, \out_fifo[0][0] [3]);
  or g41684 (n_20490, wc807, n_13893);
  not gc807 (wc807, \out_fifo[7][1] [7]);
  or g41685 (n_19686, wc808, n_13899);
  not gc808 (wc808, \out_fifo[4][0] [3]);
  or g41686 (n_19827, wc809, n_13878);
  not gc809 (wc809, \out_fifo[5][0] [4]);
  or g41687 (n_19833, wc810, n_13881);
  not gc810 (wc810, \out_fifo[2][0] [4]);
  or g41688 (n_17263, wc811, n_14702);
  not gc811 (wc811, \out_fifo[7][1] [7]);
  or g41689 (n_17264, wc812, n_14700);
  not gc812 (wc812, \out_fifo[5][1] [7]);
  or g41690 (n_17265, wc813, n_14699);
  not gc813 (wc813, \out_fifo[1][1] [7]);
  or g41691 (n_17267, wc814, n_14694);
  not gc814 (wc814, \out_fifo[6][1] [7]);
  or g41692 (n_17268, wc815, n_14695);
  not gc815 (wc815, \out_fifo[4][1] [7]);
  or g41693 (n_17269, wc816, n_14696);
  not gc816 (wc816, \out_fifo[2][1] [7]);
  or g41694 (n_15867, n_15866, wc817);
  not gc817 (wc817, n_14103);
  or g41695 (n_17270, wc818, n_14697);
  not gc818 (wc818, \out_fifo[0][1] [7]);
  or g41696 (n_17310, wc819, n_14701);
  not gc819 (wc819, \out_fifo[3][0] [5]);
  or g41697 (n_17311, wc820, n_14702);
  not gc820 (wc820, \out_fifo[7][0] [5]);
  or g41698 (n_17312, wc821, n_14700);
  not gc821 (wc821, \out_fifo[5][0] [5]);
  or g41699 (n_17313, wc822, n_14699);
  not gc822 (wc822, \out_fifo[1][0] [5]);
  or g41700 (n_18098, \data_stack_mem[3] [1], wc823);
  not gc823 (wc823, n_13926);
  or g41701 (n_17315, wc824, n_14694);
  not gc824 (wc824, \out_fifo[6][0] [5]);
  or g41702 (n_17316, wc825, n_14695);
  not gc825 (wc825, \out_fifo[4][0] [5]);
  or g41703 (n_17317, wc826, n_14696);
  not gc826 (wc826, \out_fifo[2][0] [5]);
  or g41704 (n_17318, wc827, n_14697);
  not gc827 (wc827, \out_fifo[0][0] [5]);
  or g41705 (n_17358, wc828, n_14701);
  not gc828 (wc828, \out_fifo[3][1] [5]);
  or g41706 (n_17359, wc829, n_14702);
  not gc829 (wc829, \out_fifo[7][1] [5]);
  or g41707 (n_17360, wc830, n_14700);
  not gc830 (wc830, \out_fifo[5][1] [5]);
  or g41708 (n_17361, wc831, n_14699);
  not gc831 (wc831, \out_fifo[1][1] [5]);
  or g41709 (n_20487, wc832, n_13893);
  not gc832 (wc832, \out_fifo[7][1] [5]);
  or g41710 (n_16158, wc833, n_14152);
  not gc833 (wc833, n_15497);
  or g41711 (n_17363, wc834, n_14694);
  not gc834 (wc834, \out_fifo[6][1] [5]);
  or g41712 (n_20733, wc835, n_13890);
  not gc835 (wc835, \out_fifo[3][0] [0]);
  or g41713 (n_17364, wc836, n_14695);
  not gc836 (wc836, \out_fifo[4][1] [5]);
  or g41714 (n_17365, wc837, n_14696);
  not gc837 (wc837, \out_fifo[2][1] [5]);
  or g41715 (n_17366, wc838, n_14697);
  not gc838 (wc838, \out_fifo[0][1] [5]);
  or g41716 (n_17406, wc839, n_14701);
  not gc839 (wc839, \out_fifo[3][0] [4]);
  or g41717 (n_17407, wc840, n_14702);
  not gc840 (wc840, \out_fifo[7][0] [4]);
  or g41718 (n_17408, wc841, n_14700);
  not gc841 (wc841, \out_fifo[5][0] [4]);
  or g41719 (n_17409, wc842, n_14699);
  not gc842 (wc842, \out_fifo[1][0] [4]);
  or g41720 (n_15908, n_15907, wc843);
  not gc843 (wc843, n_14236);
  or g41721 (n_19839, wc844, n_13884);
  not gc844 (wc844, \out_fifo[1][0] [4]);
  or g41722 (n_17411, wc845, n_14694);
  not gc845 (wc845, \out_fifo[6][0] [4]);
  or g41723 (n_17412, wc846, n_14695);
  not gc846 (wc846, \out_fifo[4][0] [4]);
  or g41724 (n_17413, wc847, n_14696);
  not gc847 (wc847, \out_fifo[2][0] [4]);
  or g41725 (n_17414, wc848, n_14697);
  not gc848 (wc848, \out_fifo[0][0] [4]);
  or g41726 (n_17454, wc849, n_14701);
  not gc849 (wc849, \out_fifo[3][0] [3]);
  or g41727 (n_17455, wc850, n_14702);
  not gc850 (wc850, \out_fifo[7][0] [3]);
  or g41728 (n_16056, wc851, n_14284);
  not gc851 (wc851, n_15516);
  or g41729 (n_20727, wc852, n_13887);
  not gc852 (wc852, \out_fifo[6][0] [0]);
  or g41730 (n_20721, wc853, n_13884);
  not gc853 (wc853, \out_fifo[1][0] [0]);
  or g41731 (n_17456, wc854, n_14700);
  not gc854 (wc854, \out_fifo[5][0] [3]);
  or g41732 (n_17457, wc855, n_14699);
  not gc855 (wc855, \out_fifo[1][0] [3]);
  or g41733 (n_19845, wc856, n_13887);
  not gc856 (wc856, \out_fifo[6][0] [4]);
  or g41734 (n_17459, wc857, n_14694);
  not gc857 (wc857, \out_fifo[6][0] [3]);
  or g41735 (n_17460, wc858, n_14695);
  not gc858 (wc858, \out_fifo[4][0] [3]);
  or g41736 (n_20715, wc859, n_13881);
  not gc859 (wc859, \out_fifo[2][0] [0]);
  or g41737 (n_20709, wc860, n_13878);
  not gc860 (wc860, \out_fifo[5][0] [0]);
  or g41738 (n_20703, wc861, n_13899);
  not gc861 (wc861, \out_fifo[4][1] [3]);
  or g41739 (n_20697, wc862, n_13896);
  not gc862 (wc862, \out_fifo[0][1] [3]);
  or g41740 (n_20691, wc863, n_13893);
  not gc863 (wc863, \out_fifo[7][1] [3]);
  or g41741 (n_20685, wc864, n_13890);
  not gc864 (wc864, \out_fifo[3][1] [3]);
  or g41742 (n_20679, wc865, n_13887);
  not gc865 (wc865, \out_fifo[6][1] [3]);
  or g41743 (n_20673, wc866, n_13884);
  not gc866 (wc866, \out_fifo[1][1] [3]);
  or g41744 (n_20667, wc867, n_13881);
  not gc867 (wc867, \out_fifo[2][1] [3]);
  or g41745 (n_20661, wc868, n_13878);
  not gc868 (wc868, \out_fifo[5][1] [3]);
  or g41746 (n_20646, wc869, n_13899);
  not gc869 (wc869, \out_fifo[4][1] [4]);
  or g41747 (n_20640, wc870, n_13896);
  not gc870 (wc870, \out_fifo[0][1] [4]);
  or g41748 (n_20634, wc871, n_13893);
  not gc871 (wc871, \out_fifo[7][1] [4]);
  or g41749 (n_20628, wc872, n_13890);
  not gc872 (wc872, \out_fifo[3][1] [4]);
  or g41750 (n_20622, wc873, n_13887);
  not gc873 (wc873, \out_fifo[6][1] [4]);
  or g41751 (n_20616, wc874, n_13884);
  not gc874 (wc874, \out_fifo[1][1] [4]);
  or g41752 (n_20610, wc875, n_13881);
  not gc875 (wc875, \out_fifo[2][1] [4]);
  or g41753 (n_20604, wc876, n_13878);
  not gc876 (wc876, \out_fifo[5][1] [4]);
  or g41754 (n_20598, wc877, n_13899);
  not gc877 (wc877, \out_fifo[4][1] [2]);
  or g41755 (n_20592, wc878, n_13896);
  not gc878 (wc878, \out_fifo[0][1] [2]);
  or g41756 (n_20586, wc879, n_13893);
  not gc879 (wc879, \out_fifo[7][1] [2]);
  or g41757 (n_20580, wc880, n_13890);
  not gc880 (wc880, \out_fifo[3][1] [2]);
  or g41758 (n_20574, wc881, n_13887);
  not gc881 (wc881, \out_fifo[6][1] [2]);
  or g41759 (n_20568, wc882, n_13884);
  not gc882 (wc882, \out_fifo[1][1] [2]);
  or g41760 (n_17461, wc883, n_14696);
  not gc883 (wc883, \out_fifo[2][0] [3]);
  or g41761 (n_20562, wc884, n_13881);
  not gc884 (wc884, \out_fifo[2][1] [2]);
  or g41762 (n_17462, wc885, n_14697);
  not gc885 (wc885, \out_fifo[0][0] [3]);
  or g41763 (n_17502, wc886, n_14701);
  not gc886 (wc886, \out_fifo[3][1] [4]);
  or g41764 (n_17503, wc887, n_14702);
  not gc887 (wc887, \out_fifo[7][1] [4]);
  or g41765 (n_17504, wc888, n_14700);
  not gc888 (wc888, \out_fifo[5][1] [4]);
  or g41766 (n_17505, wc889, n_14699);
  not gc889 (wc889, \out_fifo[1][1] [4]);
  or g41767 (n_19851, wc890, n_13890);
  not gc890 (wc890, \out_fifo[3][0] [4]);
  or g41768 (n_17507, wc891, n_14694);
  not gc891 (wc891, \out_fifo[6][1] [4]);
  or g41769 (n_17508, wc892, n_14695);
  not gc892 (wc892, \out_fifo[4][1] [4]);
  or g41770 (n_17509, wc893, n_14696);
  not gc893 (wc893, \out_fifo[2][1] [4]);
  or g41771 (n_17510, wc894, n_14697);
  not gc894 (wc894, \out_fifo[0][1] [4]);
  or g41772 (n_17550, wc895, n_14701);
  not gc895 (wc895, \out_fifo[3][1] [1]);
  or g41773 (n_17551, wc896, n_14702);
  not gc896 (wc896, \out_fifo[7][1] [1]);
  or g41774 (n_17552, wc897, n_14700);
  not gc897 (wc897, \out_fifo[5][1] [1]);
  or g41775 (n_17553, wc898, n_14699);
  not gc898 (wc898, \out_fifo[1][1] [1]);
  or g41776 (n_20343, wc899, n_13878);
  not gc899 (wc899, \out_fifo[5][1] [1]);
  or g41777 (n_17555, wc900, n_14694);
  not gc900 (wc900, \out_fifo[6][1] [1]);
  or g41778 (n_17556, wc901, n_14695);
  not gc901 (wc901, \out_fifo[4][1] [1]);
  nand g41779 (n_22010, n_14327, n_14333);
  or g41780 (n_22011, n_14327, n_14333);
  nand g41781 (n_14334, n_22010, n_22011);
  or g41782 (n_14141, wc902, n_15753);
  not gc902 (wc902, n_14107);
  or g41783 (n_20484, wc903, n_13893);
  not gc903 (wc903, \out_fifo[7][1] [8]);
  or g41784 (n_20481, wc904, n_13881);
  not gc904 (wc904, \out_fifo[2][1] [5]);
  or g41785 (n_16368, wc905, n_13972);
  not gc905 (wc905, n_13970);
  or g41786 (n_20442, wc906, n_13896);
  not gc906 (wc906, \out_fifo[0][1] [5]);
  or g41787 (n_16367, n_13970, n_13971);
  or g41788 (n_20460, wc907, n_13899);
  not gc907 (wc907, \out_fifo[4][1] [5]);
  or g41789 (n_20439, wc908, n_13896);
  not gc908 (wc908, \out_fifo[0][1] [6]);
  nand g41790 (n_13979, n_16322, n_16323);
  or g41791 (n_17557, wc909, n_14696);
  not gc909 (wc909, \out_fifo[2][1] [1]);
  or g41792 (n_17558, wc910, n_14697);
  not gc910 (wc910, \out_fifo[0][1] [1]);
  or g41793 (n_17598, wc911, n_14701);
  not gc911 (wc911, \out_fifo[3][0] [1]);
  or g41794 (n_17599, wc912, n_14702);
  not gc912 (wc912, \out_fifo[7][0] [1]);
  or g41795 (n_20391, wc913, n_13890);
  not gc913 (wc913, \out_fifo[3][1] [1]);
  or g41796 (n_17600, wc914, n_14700);
  not gc914 (wc914, \out_fifo[5][0] [1]);
  or g41797 (n_20457, wc915, n_13878);
  not gc915 (wc915, \out_fifo[5][1] [7]);
  or g41798 (n_17601, wc916, n_14699);
  not gc916 (wc916, \out_fifo[1][0] [1]);
  or g41799 (n_20436, wc917, n_13896);
  not gc917 (wc917, \out_fifo[0][1] [8]);
  or g41800 (n_17603, wc918, n_14694);
  not gc918 (wc918, \out_fifo[6][0] [1]);
  or g41801 (n_17604, wc919, n_14695);
  not gc919 (wc919, \out_fifo[4][0] [1]);
  or g41802 (n_17605, wc920, n_14696);
  not gc920 (wc920, \out_fifo[2][0] [1]);
  or g41803 (n_17606, wc921, n_14697);
  not gc921 (wc921, \out_fifo[0][0] [1]);
  or g41804 (n_17646, wc922, n_14701);
  not gc922 (wc922, \out_fifo[3][1] [0]);
  or g41805 (n_20556, wc923, n_13878);
  not gc923 (wc923, \out_fifo[5][1] [2]);
  or g41806 (n_20529, wc924, n_13890);
  not gc924 (wc924, \out_fifo[3][1] [8]);
  or g41807 (n_20526, wc925, n_13890);
  not gc925 (wc925, \out_fifo[3][1] [6]);
  or g41808 (n_17647, wc926, n_14702);
  not gc926 (wc926, \out_fifo[7][1] [0]);
  or g41809 (n_20523, wc927, n_13890);
  not gc927 (wc927, \out_fifo[3][1] [7]);
  or g41810 (n_20520, wc928, n_13890);
  not gc928 (wc928, \out_fifo[3][1] [5]);
  or g41811 (n_20517, wc929, n_13887);
  not gc929 (wc929, \out_fifo[6][1] [8]);
  or g41812 (n_20514, wc930, n_13887);
  not gc930 (wc930, \out_fifo[6][1] [5]);
  or g41813 (n_17648, wc931, n_14700);
  not gc931 (wc931, \out_fifo[5][1] [0]);
  or g41814 (n_17649, wc932, n_14699);
  not gc932 (wc932, \out_fifo[1][1] [0]);
  or g41815 (n_19857, wc933, n_13893);
  not gc933 (wc933, \out_fifo[7][0] [4]);
  or g41816 (n_17651, wc934, n_14694);
  not gc934 (wc934, \out_fifo[6][1] [0]);
  or g41817 (n_17652, wc935, n_14695);
  not gc935 (wc935, \out_fifo[4][1] [0]);
  or g41818 (n_17653, wc936, n_14696);
  not gc936 (wc936, \out_fifo[2][1] [0]);
  or g41819 (n_17654, wc937, n_14697);
  not gc937 (wc937, \out_fifo[0][1] [0]);
  or g41820 (n_17694, wc938, n_14701);
  not gc938 (wc938, \out_fifo[3][1] [3]);
  or g41821 (n_17695, wc939, n_14702);
  not gc939 (wc939, \out_fifo[7][1] [3]);
  or g41822 (n_17696, wc940, n_14700);
  not gc940 (wc940, \out_fifo[5][1] [3]);
  or g41823 (n_17697, wc941, n_14699);
  not gc941 (wc941, \out_fifo[1][1] [3]);
  nand g41824 (n_22012, n_14123, n_14129);
  or g41825 (n_22013, n_14123, n_14129);
  nand g41826 (n_14130, n_22012, n_22013);
  or g41827 (n_19863, wc942, n_13896);
  not gc942 (wc942, \out_fifo[0][0] [4]);
  or g41828 (n_20433, wc943, n_13899);
  not gc943 (wc943, \out_fifo[4][0] [8]);
  or g41829 (n_19869, wc944, n_13899);
  not gc944 (wc944, \out_fifo[4][0] [4]);
  nand g41830 (n_14026, n_16220, n_16221);
  or g41831 (n_20397, wc945, n_13890);
  not gc945 (wc945, \out_fifo[3][0] [8]);
  or g41832 (n_20427, wc946, n_13899);
  not gc946 (wc946, \out_fifo[4][1] [1]);
  or g41833 (n_20421, wc947, n_13896);
  not gc947 (wc947, \out_fifo[0][0] [8]);
  or g41834 (n_20403, wc948, n_13893);
  not gc948 (wc948, \out_fifo[7][1] [1]);
  or g41835 (n_20010, wc949, n_13878);
  not gc949 (wc949, \out_fifo[5][0] [5]);
  or g41836 (n_20016, wc950, n_13881);
  not gc950 (wc950, \out_fifo[2][0] [5]);
  or g41837 (n_15460, n_16386, wc951);
  not gc951 (wc951, n_13840);
  or g41838 (n_17699, wc952, n_14694);
  not gc952 (wc952, \out_fifo[6][1] [3]);
  or g41839 (n_17700, wc953, n_14695);
  not gc953 (wc953, \out_fifo[4][1] [3]);
  or g41840 (n_17701, wc954, n_14696);
  not gc954 (wc954, \out_fifo[2][1] [3]);
  or g41841 (n_17702, wc955, n_14697);
  not gc955 (wc955, \out_fifo[0][1] [3]);
  or g41842 (n_17742, wc956, n_14701);
  not gc956 (wc956, \out_fifo[3][2] [0]);
  or g41843 (n_17743, wc957, n_14702);
  not gc957 (wc957, \out_fifo[7][2] [0]);
  or g41844 (n_20022, wc958, n_13884);
  not gc958 (wc958, \out_fifo[1][0] [5]);
  or g41845 (n_17744, wc959, n_14700);
  not gc959 (wc959, \out_fifo[5][2] [0]);
  or g41846 (n_17745, wc960, n_14699);
  not gc960 (wc960, \out_fifo[1][2] [0]);
  or g41847 (n_20028, wc961, n_13887);
  not gc961 (wc961, \out_fifo[6][0] [5]);
  or g41848 (n_17747, wc962, n_14694);
  not gc962 (wc962, \out_fifo[6][2] [0]);
  or g41849 (n_17748, wc963, n_14695);
  not gc963 (wc963, \out_fifo[4][2] [0]);
  or g41850 (n_20034, wc964, n_13890);
  not gc964 (wc964, \out_fifo[3][0] [5]);
  or g41851 (n_17749, wc965, n_14696);
  not gc965 (wc965, \out_fifo[2][2] [0]);
  or g41852 (n_17750, wc966, n_14697);
  not gc966 (wc966, \out_fifo[0][2] [0]);
  or g41853 (n_17790, wc967, n_14696);
  not gc967 (wc967, \out_fifo[2][0] [6]);
  or g41854 (n_17791, wc968, n_14695);
  not gc968 (wc968, \out_fifo[4][0] [6]);
  or g41855 (n_20040, wc969, n_13893);
  not gc969 (wc969, \out_fifo[7][0] [5]);
  or g41856 (n_17792, wc970, n_14694);
  not gc970 (wc970, \out_fifo[6][0] [6]);
  or g41857 (n_17793, wc971, n_14697);
  not gc971 (wc971, \out_fifo[0][0] [6]);
  or g41858 (n_20046, wc972, n_13896);
  not gc972 (wc972, \out_fifo[0][0] [5]);
  or g41859 (n_20052, wc973, n_13899);
  not gc973 (wc973, \out_fifo[4][0] [5]);
  or g41860 (n_17795, wc974, n_14699);
  not gc974 (wc974, \out_fifo[1][0] [6]);
  or g41861 (n_17796, wc975, n_14700);
  not gc975 (wc975, \out_fifo[5][0] [6]);
  or g41862 (n_17797, wc976, n_14701);
  not gc976 (wc976, \out_fifo[3][0] [6]);
  or g41863 (n_14109, wc977, n_15741);
  not gc977 (wc977, n_14107);
  or g41864 (n_20109, wc978, n_13878);
  not gc978 (wc978, \out_fifo[5][0] [6]);
  or g41865 (n_20115, wc979, n_13881);
  not gc979 (wc979, \out_fifo[2][0] [6]);
  or g41866 (n_20121, wc980, n_13884);
  not gc980 (wc980, \out_fifo[1][0] [6]);
  or g41867 (n_20127, wc981, n_13887);
  not gc981 (wc981, \out_fifo[6][0] [6]);
  or g41868 (n_20133, wc982, n_13890);
  not gc982 (wc982, \out_fifo[3][0] [6]);
  nand g41869 (n_22014, n_14274, n_14280);
  or g41870 (n_22015, n_14274, n_14280);
  nand g41871 (n_14281, n_22014, n_22015);
  or g41872 (n_20139, wc983, n_13893);
  not gc983 (wc983, \out_fifo[7][0] [6]);
  or g41873 (n_20415, wc984, n_13896);
  not gc984 (wc984, \out_fifo[0][1] [1]);
  or g41874 (n_20145, wc985, n_13896);
  not gc985 (wc985, \out_fifo[0][0] [6]);
  or g41875 (n_20151, wc986, n_13899);
  not gc986 (wc986, \out_fifo[4][0] [6]);
  nand g41876 (n_22016, n_13965, n_14004);
  or g41877 (n_22017, n_13965, n_14004);
  nand g41878 (n_14005, n_22016, n_22017);
  or g41879 (n_20409, wc987, n_13893);
  not gc987 (wc987, \out_fifo[7][0] [8]);
  or g41880 (n_17798, wc988, n_14702);
  not gc988 (wc988, \out_fifo[7][0] [6]);
  or g41883 (n_17838, wc989, n_14696);
  not gc989 (wc989, \out_fifo[2][0] [2]);
  or g41884 (n_16434, wc990, n_13926);
  not gc990 (wc990, n_13914);
  or g41885 (n_17839, wc991, n_14695);
  not gc991 (wc991, \out_fifo[4][0] [2]);
  or g41886 (n_17840, wc992, n_14694);
  not gc992 (wc992, \out_fifo[6][0] [2]);
  or g41887 (n_20373, wc993, n_13884);
  not gc993 (wc993, \out_fifo[1][0] [8]);
  or g41888 (n_17841, wc994, n_14697);
  not gc994 (wc994, \out_fifo[0][0] [2]);
  or g41889 (n_20454, wc995, n_13878);
  not gc995 (wc995, \out_fifo[5][1] [5]);
  or g41890 (n_20451, wc996, n_13878);
  not gc996 (wc996, \out_fifo[5][1] [6]);
  or g41891 (n_20379, wc997, n_13887);
  not gc997 (wc997, \out_fifo[6][1] [1]);
  or g41892 (n_17843, wc998, n_14699);
  not gc998 (wc998, \out_fifo[1][0] [2]);
  or g41893 (n_17844, wc999, n_14700);
  not gc999 (wc999, \out_fifo[5][0] [2]);
  or g41894 (n_17845, wc1000, n_14701);
  not gc1000 (wc1000, \out_fifo[3][0] [2]);
  or g41895 (n_17846, wc1001, n_14702);
  not gc1001 (wc1001, \out_fifo[7][0] [2]);
  or g41896 (n_17886, wc1002, n_14696);
  not gc1002 (wc1002, \out_fifo[2][2] [8]);
  or g41897 (n_17887, wc1003, n_14695);
  not gc1003 (wc1003, \out_fifo[4][2] [8]);
  or g41898 (n_17888, wc1004, n_14694);
  not gc1004 (wc1004, \out_fifo[6][2] [8]);
  or g41899 (n_17889, wc1005, n_14697);
  not gc1005 (wc1005, \out_fifo[0][2] [8]);
  nand g41900 (n_14682, n_16100, n_16101);
  or g41901 (n_20448, wc1006, n_13878);
  not gc1006 (wc1006, \out_fifo[5][1] [8]);
  or g41902 (n_17891, wc1007, n_14699);
  not gc1007 (wc1007, \out_fifo[1][2] [8]);
  or g41903 (n_17892, wc1008, n_14700);
  not gc1008 (wc1008, \out_fifo[5][2] [8]);
  or g41904 (n_17893, wc1009, n_14701);
  not gc1009 (wc1009, \out_fifo[3][2] [8]);
  or g41905 (n_17894, wc1010, n_14702);
  not gc1010 (wc1010, \out_fifo[7][2] [8]);
  or g41906 (n_17934, wc1011, n_14696);
  not gc1011 (wc1011, \out_fifo[2][2] [1]);
  or g41907 (n_17935, wc1012, n_14695);
  not gc1012 (wc1012, \out_fifo[4][2] [1]);
  or g41908 (n_17936, wc1013, n_14694);
  not gc1013 (wc1013, \out_fifo[6][2] [1]);
  or g41909 (n_17937, wc1014, n_14697);
  not gc1014 (wc1014, \out_fifo[0][2] [1]);
  or g41910 (n_20445, wc1015, n_13896);
  not gc1015 (wc1015, \out_fifo[0][1] [7]);
  or g41911 (n_17939, wc1016, n_14699);
  not gc1016 (wc1016, \out_fifo[1][2] [1]);
  or g41912 (n_20208, wc1017, n_13878);
  not gc1017 (wc1017, \out_fifo[5][0] [7]);
  or g41913 (n_17940, wc1018, n_14700);
  not gc1018 (wc1018, \out_fifo[5][2] [1]);
  or g41914 (n_17941, wc1019, n_14701);
  not gc1019 (wc1019, \out_fifo[3][2] [1]);
  nand g41915 (n_14262, n_15717, n_20829);
  or g41916 (n_17942, wc1020, n_14702);
  not gc1020 (wc1020, \out_fifo[7][2] [1]);
  or g41917 (n_17982, wc1021, n_14696);
  not gc1021 (wc1021, \out_fifo[2][1] [2]);
  or g41918 (n_17983, wc1022, n_14695);
  not gc1022 (wc1022, \out_fifo[4][1] [2]);
  or g41919 (n_17984, wc1023, n_14694);
  not gc1023 (wc1023, \out_fifo[6][1] [2]);
  or g41920 (n_17985, wc1024, n_14697);
  not gc1024 (wc1024, \out_fifo[0][1] [2]);
  or g41921 (n_20511, wc1025, n_13887);
  not gc1025 (wc1025, \out_fifo[6][1] [7]);
  or g41922 (n_17987, wc1026, n_14699);
  not gc1026 (wc1026, \out_fifo[1][1] [2]);
  or g41923 (n_17988, wc1027, n_14700);
  not gc1027 (wc1027, \out_fifo[5][1] [2]);
  or g41924 (n_17989, wc1028, n_14701);
  not gc1028 (wc1028, \out_fifo[3][1] [2]);
  nand g41925 (n_14679, n_16271, n_16272);
  nand g41926 (n_16280, n_15463, data_stack_pointer[3]);
  or g41927 (n_17990, wc1029, n_14702);
  not gc1029 (wc1029, \out_fifo[7][1] [2]);
  or g41928 (n_18030, wc1030, n_14696);
  not gc1030 (wc1030, \out_fifo[2][2] [9]);
  or g41929 (n_18031, wc1031, n_14695);
  not gc1031 (wc1031, \out_fifo[4][2] [9]);
  or g41930 (n_20214, wc1032, n_13881);
  not gc1032 (wc1032, \out_fifo[2][0] [7]);
  or g41931 (n_20508, wc1033, n_13887);
  not gc1033 (wc1033, \out_fifo[6][1] [6]);
  or g41932 (n_20220, wc1034, n_13884);
  not gc1034 (wc1034, \out_fifo[1][0] [7]);
  or g41933 (n_20505, wc1035, n_13884);
  not gc1035 (wc1035, \out_fifo[1][1] [5]);
  or g41934 (n_16362, wc1036, n_13972);
  not gc1036 (wc1036, n_13926);
  or g41935 (n_16361, n_13926, n_13971);
  nand g41936 (n_13989, n_16328, n_16329);
  or g41937 (n_20385, wc1037, n_13887);
  not gc1037 (wc1037, \out_fifo[6][0] [8]);
  or g41938 (n_20349, wc1038, n_13878);
  not gc1038 (wc1038, \out_fifo[5][0] [8]);
  or g41939 (n_18032, wc1039, n_14694);
  not gc1039 (wc1039, \out_fifo[6][2] [9]);
  or g41940 (n_18033, wc1040, n_14697);
  not gc1040 (wc1040, \out_fifo[0][2] [9]);
  or g41941 (n_20478, wc1041, n_13881);
  not gc1041 (wc1041, \out_fifo[2][1] [6]);
  nand g41942 (n_14063, n_16214, n_16215);
  or g41943 (n_20475, wc1042, n_13881);
  not gc1042 (wc1042, \out_fifo[2][1] [7]);
  or g41944 (n_13857, n_13856, wc1043);
  not gc1043 (wc1043, n_16443);
  or g41945 (n_20355, wc1044, n_13881);
  not gc1044 (wc1044, \out_fifo[2][1] [1]);
  or g41946 (n_14610, n_14587, wc1045);
  not gc1045 (wc1045, n_16446);
  or g41947 (n_20472, wc1046, n_13881);
  not gc1046 (wc1046, \out_fifo[2][1] [8]);
  or g41948 (n_18035, wc1047, n_14699);
  not gc1047 (wc1047, \out_fifo[1][2] [9]);
  nand g41949 (n_14684, n_16451, n_16452);
  or g41950 (n_18036, wc1048, n_14700);
  not gc1048 (wc1048, \out_fifo[5][2] [9]);
  or g41951 (n_18037, wc1049, n_14701);
  not gc1049 (wc1049, \out_fifo[3][2] [9]);
  or g41952 (n_14588, n_14587, wc1050);
  not gc1050 (wc1050, n_16455);
  or g41953 (n_18038, wc1051, n_14702);
  not gc1051 (wc1051, \out_fifo[7][2] [9]);
  or g41954 (n_14630, n_13856, wc1052);
  not gc1052 (wc1052, n_16458);
  or g41955 (n_18078, wc1053, n_14696);
  not gc1053 (wc1053, \out_fifo[2][1] [8]);
  or g41956 (n_14598, n_14587, wc1054);
  not gc1054 (wc1054, n_16461);
  or g41957 (n_18079, wc1055, n_14695);
  not gc1055 (wc1055, \out_fifo[4][1] [8]);
  or g41958 (n_14620, n_14587, wc1056);
  not gc1056 (wc1056, n_16464);
  or g41959 (n_18104, wc1057, n_13970);
  not gc1057 (wc1057, \data_stack_mem[3] [1]);
  or g41960 (n_14640, n_13856, wc1058);
  not gc1058 (wc1058, n_16467);
  or g41961 (n_18080, wc1059, n_14694);
  not gc1059 (wc1059, \out_fifo[6][1] [8]);
  or g41962 (n_18081, wc1060, n_14697);
  not gc1060 (wc1060, \out_fifo[0][1] [8]);
  or g41963 (n_13859, data_stack_pointer[2], n_20805);
  or g41964 (n_16520, n_13879, n_13876);
  or g41965 (n_16521, wc1061, n_13878);
  not gc1061 (wc1061, \out_fifo[5][2] [8]);
  or g41966 (n_16526, n_13882, n_13876);
  or g41967 (n_20469, wc1062, n_13899);
  not gc1062 (wc1062, \out_fifo[4][1] [7]);
  or g41968 (n_16527, wc1063, n_13881);
  not gc1063 (wc1063, \out_fifo[2][2] [8]);
  or g41969 (n_16532, n_13885, n_13876);
  or g41970 (n_18083, wc1064, n_14699);
  not gc1064 (wc1064, \out_fifo[1][1] [8]);
  or g41971 (n_16533, wc1065, n_13884);
  not gc1065 (wc1065, \out_fifo[1][2] [8]);
  or g41972 (n_16538, n_13888, n_13876);
  or g41973 (n_16539, wc1066, n_13887);
  not gc1066 (wc1066, \out_fifo[6][2] [8]);
  or g41974 (n_16544, n_13891, n_13876);
  or g41975 (n_16545, wc1067, n_13890);
  not gc1067 (wc1067, \out_fifo[3][2] [8]);
  or g41976 (n_16550, n_13894, n_13876);
  nand g41977 (n_14245, n_15621, n_20814);
  or g41978 (n_18084, wc1068, n_14700);
  not gc1068 (wc1068, \out_fifo[5][1] [8]);
  or g41979 (n_18085, wc1069, n_14701);
  not gc1069 (wc1069, \out_fifo[3][1] [8]);
  or g41980 (n_18086, wc1070, n_14702);
  not gc1070 (wc1070, \out_fifo[7][1] [8]);
  or g41981 (n_19242, wc1071, n_13878);
  not gc1071 (wc1071, \out_fifo[5][0] [1]);
  or g41982 (n_19248, wc1072, n_13881);
  not gc1072 (wc1072, \out_fifo[2][0] [1]);
  or g41983 (n_19254, wc1073, n_13884);
  not gc1073 (wc1073, \out_fifo[1][0] [1]);
  or g41984 (n_16551, wc1074, n_13893);
  not gc1074 (wc1074, \out_fifo[7][2] [8]);
  or g41985 (n_16556, n_13897, n_13876);
  or g41986 (n_16557, wc1075, n_13896);
  not gc1075 (wc1075, \out_fifo[0][2] [8]);
  or g41987 (n_16562, n_13900, n_13876);
  or g41988 (n_16563, wc1076, n_13899);
  not gc1076 (wc1076, \out_fifo[4][2] [8]);
  or g41989 (n_16568, wc1077, n_14584);
  not gc1077 (wc1077, sh_reg_in[4]);
  or g41990 (n_16574, wc1078, n_14584);
  not gc1078 (wc1078, sh_reg_in[5]);
  or g41991 (n_16580, wc1079, n_14584);
  not gc1079 (wc1079, sh_reg_in[6]);
  or g41992 (n_16586, wc1080, n_14584);
  not gc1080 (wc1080, sh_reg_in[3]);
  or g41993 (n_16592, wc1081, n_14584);
  not gc1081 (wc1081, sh_reg_in[2]);
  or g41994 (n_16598, wc1082, n_14584);
  not gc1082 (wc1082, sh_reg_in[1]);
  or g41995 (n_16604, wc1083, n_14584);
  not gc1083 (wc1083, sh_reg_in[0]);
  nand g41996 (n_16433, n_14980, n_13925);
  or g41997 (n_13900, n_13837, wc1084);
  not gc1084 (wc1084, rst_n);
  nand g41998 (n_13899, rst_n, n_13837);
  or g41999 (n_13897, n_13846, wc1085);
  not gc1085 (wc1085, rst_n);
  nand g42000 (n_13896, rst_n, n_13846);
  or g42001 (n_15907, n_15906, wc1086);
  not gc1086 (wc1086, n_14241);
  or g42002 (n_13894, n_13830, wc1087);
  not gc1087 (wc1087, rst_n);
  nand g42003 (n_13893, rst_n, n_13830);
  or g42004 (n_16322, wc1088, n_13978);
  not gc1088 (wc1088, n_15310);
  or g42005 (n_14284, n_15726, wc1089);
  not gc1089 (wc1089, \data_stack_mem[0] [5]);
  nand g42006 (n_22019, n_14369, n_14466);
  or g42007 (n_22020, n_14369, n_14466);
  nand g42008 (n_14467, n_22019, n_22020);
  or g42009 (n_16323, n_15310, wc1090);
  not gc1090 (wc1090, n_13978);
  or g42010 (n_16328, wc1091, n_13988);
  not gc1091 (wc1091, n_15372);
  or g42011 (n_16329, n_15372, wc1092);
  not gc1092 (wc1092, n_13988);
  or g42012 (n_15866, n_15865, wc1093);
  not gc1093 (wc1093, n_14102);
  nand g42013 (n_22021, n_13998, n_14003);
  or g42014 (n_22022, n_13998, n_14003);
  nand g42015 (n_14004, n_22021, n_22022);
  nand g42016 (n_22023, n_14328, n_14332);
  or g42017 (n_22024, n_14328, n_14332);
  nand g42018 (n_14333, n_22023, n_22024);
  or g42019 (n_15845, n_15844, wc1094);
  not gc1094 (wc1094, n_14021);
  or g42020 (n_13891, n_13840, wc1095);
  not gc1095 (wc1095, rst_n);
  nand g42021 (n_16220, n_15340, n_13924);
  or g42022 (n_14584, n_13869, n_14583);
  nand g42023 (n_13890, rst_n, n_13840);
  or g42024 (n_13888, n_13833, wc1096);
  not gc1096 (wc1096, rst_n);
  or g42025 (n_14641, n_13858, n_13869);
  nand g42026 (n_13887, rst_n, n_13833);
  or g42027 (n_14699, n_13903, n_14698);
  nand g42028 (n_22025, n_14045, n_14050);
  or g42029 (n_22026, n_14045, n_14050);
  nand g42030 (n_14051, n_22025, n_22026);
  or g42031 (n_14700, n_13904, n_14698);
  or g42032 (n_16214, n_13974, wc1097);
  not gc1097 (wc1097, n_15321);
  or g42033 (n_14702, n_13902, n_14698);
  or g42034 (n_16167, n_16166, wc1098);
  not gc1098 (wc1098, n_14020);
  or g42035 (n_14701, n_13905, n_14698);
  or g42036 (n_13885, n_13844, wc1099);
  not gc1099 (wc1099, rst_n);
  nand g42037 (n_13884, rst_n, n_13844);
  or g42038 (n_14697, n_13903, n_14693);
  or g42039 (n_14694, n_13902, n_14693);
  or g42040 (n_13882, n_13842, wc1100);
  not gc1100 (wc1100, rst_n);
  or g42041 (n_14008, n_15705, wc1101);
  not gc1101 (wc1101, \data_stack_mem[0] [1]);
  or g42042 (n_16350, \data_stack_mem[2] [2], wc1102);
  not gc1102 (wc1102, n_14031);
  nand g42043 (n_13881, rst_n, n_13842);
  or g42044 (n_13879, n_13835, wc1103);
  not gc1103 (wc1103, rst_n);
  or g42045 (n_14695, n_13904, n_14693);
  or g42046 (n_14696, n_13905, n_14693);
  or g42047 (n_15887, n_15886, wc1104);
  not gc1104 (wc1104, n_14170);
  nand g42048 (n_15741, n_15739, n_15740);
  nand g42049 (n_13878, rst_n, n_13835);
  or g42050 (n_14597, n_14583, n_14987);
  nand g42051 (n_22027, n_14124, n_14128);
  or g42052 (n_22028, n_14124, n_14128);
  nand g42053 (n_14129, n_22027, n_22028);
  nand g42054 (n_16344, \data_stack_mem[2] [2], n_14065);
  or g42055 (n_14619, n_14583, n_14986);
  or g42056 (n_16046, n_16045, wc1105);
  not gc1105 (wc1105, n_14169);
  nand g42057 (n_16386, n_14909, n_16385);
  or g42058 (n_15824, n_15823, wc1106);
  not gc1106 (wc1106, n_13972);
  nand g42061 (n_15753, n_15751, n_15752);
  or g42062 (n_14355, n_15987, wc1107);
  not gc1107 (wc1107, n_14308);
  or g42063 (n_16068, n_14179, n_14176);
  or g42064 (n_16070, n_14177, wc1108);
  not gc1108 (wc1108, n_14179);
  or g42065 (n_20832, n_16317, n_13858);
  or g42066 (n_15486, wc1109, n_15648);
  not gc1109 (wc1109, n_13904);
  or g42067 (n_16081, n_14177, n_14198);
  or g42068 (n_16080, n_14176, wc1110);
  not gc1110 (wc1110, n_14198);
  nand g42069 (n_22030, n_14236, n_14279);
  or g42070 (n_22031, n_14236, n_14279);
  nand g42071 (n_14280, n_22030, n_22031);
  or g42072 (n_16101, data_stack_pointer[2], n_16099);
  nand g42073 (n_22032, n_14209, n_14212);
  or g42074 (n_22033, n_14209, n_14212);
  nand g42075 (n_14213, n_22032, n_22033);
  nand g42076 (n_14678, n_16106, n_16107);
  nand g42077 (n_20814, n_15041, n_14179);
  or g42078 (n_13950, n_13949, n_16290);
  or g42079 (n_20805, n_15552, n_13858);
  or g42080 (n_16464, n_14583, wc1111);
  not gc1111 (wc1111, n_14986);
  or g42081 (n_16461, n_14583, wc1112);
  not gc1112 (wc1112, n_14987);
  nand g42082 (n_15463, n_16148, n_16149);
  or g42083 (n_16027, n_16026, wc1113);
  not gc1113 (wc1113, n_14993);
  or g42084 (n_16455, wc1114, n_14583);
  not gc1114 (wc1114, n_13869);
  nand g42085 (n_16451, n_14651, rst_n);
  or g42086 (n_15929, n_15928, wc1115);
  not gc1115 (wc1115, n_14304);
  or g42087 (n_16446, n_14583, wc1116);
  not gc1116 (wc1116, n_14608);
  nand g42088 (n_20829, n_15442, n_14198);
  or g42089 (n_14683, n_16356, n_13855);
  or g42090 (n_16271, n_16270, wc1117);
  not gc1117 (wc1117, data_stack_pointer[0]);
  or g42091 (n_14650, n_16353, n_13855);
  or g42092 (n_14473, n_16008, wc1118);
  not gc1118 (wc1118, n_14388);
  nand g42093 (n_14587, n_16337, n_16270);
  nand g42094 (n_13856, n_16332, n_13855);
  nand g42095 (n_16272, n_15462, data_stack_pointer[1]);
  or g42096 (n_14609, n_16279, wc1119);
  not gc1119 (wc1119, data_stack_pointer[1]);
  or g42097 (n_15946, n_15945, wc1120);
  not gc1120 (wc1120, n_14376);
  or g42098 (n_14152, n_15999, wc1121);
  not gc1121 (wc1121, n_14104);
  nand g42099 (n_14750, n_13907, n_16287);
  or g42100 (n_14651, wc1122, n_13854);
  not gc1122 (wc1122, n_16317);
  nand g42101 (n_14748, n_13907, n_16284);
  nand g42102 (n_16332, n_13854, rst_n);
  or g42103 (n_16279, n_14608, n_14677);
  or g42104 (n_15945, n_15944, wc1123);
  not gc1123 (wc1123, n_14373);
  or g42105 (n_16008, n_16007, wc1124);
  not gc1124 (wc1124, n_14377);
  or g42106 (n_16353, n_13868, n_13854);
  or g42107 (n_16270, n_14586, n_14582);
  nand g42108 (n_14749, n_13907, n_16233);
  or g42109 (n_13858, n_13854, wc1125);
  not gc1125 (wc1125, rst_n);
  or g42110 (n_16356, n_14607, n_13854);
  nand g42111 (n_13909, n_13907, n_16227);
  nand g42112 (n_13908, n_13907, n_16224);
  or g42113 (n_15928, n_15927, wc1126);
  not gc1126 (wc1126, n_14298);
  nand g42114 (n_19234, \data_stack_mem[0] [0], n_13912);
  nand g42115 (n_16149, n_14680, rst_n);
  nand g42116 (n_15462, n_14866, n_16143);
  or g42117 (n_16026, n_16025, wc1127);
  not gc1127 (wc1127, n_14967);
  or g42118 (n_16106, data_stack_pointer[0], n_14677);
  or g42119 (n_16099, n_13915, n_14677);
  or g42120 (n_16100, n_13855, wc1128);
  not gc1128 (wc1128, n_14680);
  nand g42121 (n_22034, n_14275, n_14278);
  or g42122 (n_22035, n_14275, n_14278);
  nand g42123 (n_14279, n_22034, n_22035);
  or g42124 (n_13949, n_13948, n_16170);
  nand g42125 (n_22036, n_14170, n_14211);
  or g42126 (n_22037, n_14170, n_14211);
  nand g42127 (n_14212, n_22036, n_22037);
  or g42128 (n_15987, n_15986, wc1129);
  not gc1129 (wc1129, n_14305);
  nand g42129 (n_14198, n_15711, n_20826);
  nand g42130 (n_20200, \data_stack_mem[0] [6], n_13912);
  or g42131 (n_19420, wc1130, n_13876);
  not gc1130 (wc1130, \data_stack_mem[0] [1]);
  nand g42132 (n_15648, n_15646, n_15647);
  or g42133 (n_14914, n_13939, n_13937);
  nand g42138 (n_14179, n_15618, n_20811);
  nand g42139 (n_22040, out_fifo_write_pointer[1], n_13829);
  or g42140 (n_22041, out_fifo_write_pointer[1], n_13829);
  nand g42141 (n_15461, n_22040, n_22041);
  or g42142 (n_15823, n_15822, wc1131);
  not gc1131 (wc1131, n_13965);
  or g42143 (n_15751, n_15750, wc1132);
  not gc1132 (wc1132, n_13920);
  nand g42144 (n_13877, n_13870, n_13876);
  nand g42145 (n_16385, out_fifo_write_pointer[2], n_13829);
  nand g42146 (n_20002, \data_stack_mem[0] [4], n_13912);
  or g42147 (n_16045, n_16044, wc1133);
  not gc1133 (wc1133, n_14167);
  nand g42148 (n_22042, n_14100, n_14127);
  or g42149 (n_22043, n_14100, n_14127);
  nand g42150 (n_14128, n_22042, n_22043);
  or g42151 (n_15886, n_15885, wc1134);
  not gc1134 (wc1134, n_14172);
  or g42152 (n_15705, n_15704, wc1135);
  not gc1135 (wc1135, n_13975);
  or g42153 (n_15740, n_15738, wc1136);
  not gc1136 (wc1136, n_13920);
  nand g42154 (n_19636, \data_stack_mem[0] [2], n_13912);
  or g42155 (n_14065, wc1137, n_15801);
  not gc1137 (wc1137, n_14029);
  nand g42156 (n_16215, \data_stack_mem[2] [1], n_13978);
  or g42157 (n_16166, n_14075, n_16165);
  nand g42158 (n_22044, n_14021, n_14049);
  or g42159 (n_22045, n_14021, n_14049);
  nand g42160 (n_14050, n_22044, n_22045);
  or g42161 (n_14031, wc1138, n_15789);
  not gc1138 (wc1138, n_14029);
  or g42162 (n_14698, wc1139, n_13907);
  not gc1139 (wc1139, out_fifo_read_pointer[0]);
  or g42163 (n_14693, out_fifo_read_pointer[0], n_13907);
  or g42164 (n_16221, \data_stack_mem[2] [1], wc1140);
  not gc1140 (wc1140, n_13988);
  nand g42165 (n_22046, n_14304, n_14331);
  or g42166 (n_22047, n_14304, n_14331);
  nand g42167 (n_14332, n_22046, n_22047);
  or g42168 (n_15865, n_15864, wc1141);
  not gc1141 (wc1141, n_14100);
  or g42169 (n_15844, n_15843, wc1142);
  not gc1142 (wc1142, n_14015);
  nand g42170 (n_22048, n_13999, n_14002);
  or g42171 (n_22049, n_13999, n_14002);
  nand g42172 (n_14003, n_22048, n_22049);
  or g42173 (n_14583, wc1143, n_14582);
  not gc1143 (wc1143, data_stack_pointer[1]);
  nand g42174 (n_15372, n_16139, n_16140);
  or g42175 (n_15726, n_15725, wc1144);
  not gc1144 (wc1144, n_14242);
  nand g42176 (n_22050, n_14462, n_14465);
  or g42177 (n_22051, n_14462, n_14465);
  nand g42178 (n_14466, n_22050, n_22051);
  or g42179 (n_15906, n_15905, wc1145);
  not gc1145 (wc1145, n_14233);
  or g42180 (n_20098, wc1146, n_13876);
  not gc1146 (wc1146, \data_stack_mem[0] [5]);
  nand g42181 (n_15310, n_16124, n_16125);
  nand g42182 (n_19819, \data_stack_mem[0] [3], n_13912);
  nand g42183 (n_13925, n_16196, n_16197);
  or g42184 (n_15999, n_15998, wc1147);
  not gc1147 (wc1147, n_14101);
  or g42185 (n_17314, wc1148, n_13816);
  not gc1148 (wc1148, sh_reg_out[4]);
  or g42186 (n_15998, n_15997, wc1149);
  not gc1149 (wc1149, n_14099);
  or g42191 (n_17362, wc1150, n_13816);
  not gc1150 (wc1150, sh_reg_out[14]);
  or g42194 (n_15905, n_15904, wc1151);
  not gc1151 (wc1151, n_14274);
  or g42195 (n_17410, wc1152, n_13816);
  not gc1152 (wc1152, sh_reg_out[3]);
  nand g42198 (n_22056, out_fifo_read_pointer[1], n_14672);
  or g42199 (n_22057, out_fifo_read_pointer[1], n_14672);
  nand g42200 (n_15485, n_22056, n_22057);
  or g42201 (n_16025, n_16024, wc1153);
  not gc1153 (wc1153, n_14951);
  or g42202 (n_15646, n_13905, n_14672);
  nand g42203 (n_15647, out_fifo_read_pointer[2], n_14672);
  or g42204 (n_15725, n_15724, wc1154);
  not gc1154 (wc1154, n_14239);
  or g42205 (n_17458, wc1155, n_13816);
  not gc1155 (wc1155, sh_reg_out[2]);
  or g42206 (n_17506, wc1156, n_13816);
  not gc1156 (wc1156, sh_reg_out[13]);
  or g42207 (n_14582, n_14911, wc1157);
  not gc1157 (wc1157, rst_n);
  or g42208 (n_14915, n_13913, n_13940);
  or g42209 (n_15986, n_15985, wc1158);
  not gc1158 (wc1158, n_14303);
  or g42210 (n_17554, wc1159, n_13816);
  not gc1159 (wc1159, sh_reg_out[10]);
  nand g42211 (n_15789, n_15787, n_15788);
  nand g42212 (n_15443, n_13945, n_15960);
  or g42213 (n_15752, n_14106, wc1160);
  not gc1160 (wc1160, n_14140);
  nand g42214 (n_15455, n_13945, n_15966);
  or g42215 (n_15750, wc1161, n_14140);
  not gc1161 (wc1161, n_14105);
  nand g42216 (n_22058, n_14046, n_14048);
  or g42217 (n_22059, n_14046, n_14048);
  nand g42218 (n_14049, n_22058, n_22059);
  nand g42223 (n_13876, n_15518, n_13870);
  or g42224 (n_16140, wc1162, n_13973);
  not gc1162 (wc1162, n_13924);
  or g42225 (n_16139, n_13924, n_13975);
  or g42226 (n_17842, wc1163, n_13816);
  not gc1163 (wc1163, sh_reg_out[1]);
  or g42227 (n_14677, n_13853, n_14676);
  or g42228 (n_16044, n_16043, wc1164);
  not gc1164 (wc1164, n_14879);
  or g42229 (n_17602, wc1165, n_13816);
  not gc1165 (wc1165, sh_reg_out[0]);
  or g42230 (n_17650, wc1166, n_13816);
  not gc1166 (wc1166, sh_reg_out[9]);
  or g42233 (n_17890, wc1167, n_13816);
  not gc1167 (wc1167, sh_reg_out[27]);
  nand g42234 (n_22063, n_14172, n_14210);
  or g42235 (n_22064, n_14172, n_14210);
  nand g42236 (n_14211, n_22063, n_22064);
  or g42237 (n_15864, n_15863, wc1168);
  not gc1168 (wc1168, n_14094);
  or g42238 (n_17938, wc1169, n_13816);
  not gc1169 (wc1169, sh_reg_out[20]);
  nand g42239 (n_22065, n_14306, n_14330);
  or g42240 (n_22066, n_14306, n_14330);
  nand g42241 (n_14331, n_22065, n_22066);
  or g42242 (n_14680, n_13853, wc1170);
  not gc1170 (wc1170, n_16086);
  nand g42243 (n_22067, n_14102, n_14126);
  or g42244 (n_22068, n_14102, n_14126);
  nand g42245 (n_14127, n_22067, n_22068);
  or g42246 (n_13978, wc1171, n_15765);
  not gc1171 (wc1171, n_14871);
  or g42247 (n_17986, wc1172, n_13816);
  not gc1172 (wc1172, sh_reg_out[11]);
  or g42248 (n_13988, wc1173, n_15777);
  not gc1173 (wc1173, n_14871);
  nand g42249 (n_15373, n_13945, n_15954);
  or g42250 (n_16107, wc1174, n_14866);
  not gc1174 (wc1174, data_stack_pointer[0]);
  nand g42251 (n_15801, n_15799, n_15800);
  or g42252 (n_16125, n_13973, wc1175);
  not gc1175 (wc1175, n_13974);
  or g42253 (n_14629, n_14866, wc1176);
  not gc1176 (wc1176, n_16110);
  or g42254 (n_16143, data_stack_pointer[0], n_14676);
  nand g42255 (n_20826, n_15433, n_14140);
  or g42256 (n_13907, wc1177, n_13906);
  not gc1177 (wc1177, n_15459);
  or g42257 (n_16148, data_stack_pointer[2], n_14676);
  or g42258 (n_15843, n_15842, wc1178);
  not gc1178 (wc1178, n_14045);
  or g42259 (n_17698, wc1179, n_13816);
  not gc1179 (wc1179, sh_reg_out[12]);
  or g42260 (n_16224, wc1180, n_13816);
  not gc1180 (wc1180, dout_valid);
  or g42261 (n_13948, wc1181, n_16032);
  not gc1181 (wc1181, n_15510);
  or g42262 (n_16227, sh_reg_out_bit_counter[0], n_13816);
  or g42263 (n_15927, n_15926, wc1182);
  not gc1182 (wc1182, n_14306);
  nand g42264 (n_22069, n_13972, n_14001);
  or g42265 (n_22070, n_13972, n_14001);
  nand g42266 (n_14002, n_22069, n_22070);
  or g42267 (n_17746, wc1183, n_13816);
  not gc1183 (wc1183, sh_reg_out[19]);
  or g42268 (n_14075, n_15990, wc1184);
  not gc1184 (wc1184, n_14025);
  or g42269 (n_16233, n_16232, n_13816);
  nand g42270 (n_13912, n_16089, n_13910);
  or g42271 (n_17122, wc1185, n_13816);
  not gc1185 (wc1185, sh_reg_out[7]);
  nand g42272 (n_22071, n_14373, n_14464);
  or g42273 (n_22072, n_14373, n_14464);
  nand g42274 (n_14465, n_22071, n_22072);
  or g42275 (n_15704, n_15703, wc1186);
  not gc1186 (wc1186, n_13971);
  or g42276 (n_17794, wc1187, n_13816);
  not gc1187 (wc1187, sh_reg_out[5]);
  or g42277 (n_16007, n_16006, wc1188);
  not gc1188 (wc1188, n_14372);
  or g42278 (n_17170, wc1189, n_13816);
  not gc1189 (wc1189, sh_reg_out[15]);
  or g42279 (n_16284, wc1190, n_13816);
  not gc1190 (wc1190, n_15473);
  nand g42280 (n_15430, n_13945, n_15957);
  or g42285 (n_16287, wc1191, n_13816);
  not gc1191 (wc1191, n_15474);
  nand g42286 (n_15447, n_13945, n_15963);
  or g42287 (n_17218, wc1192, n_13816);
  not gc1192 (wc1192, sh_reg_out[6]);
  nand g42288 (n_15738, n_14105, n_14108);
  nand g42289 (n_15301, n_13945, n_15951);
  or g42290 (n_15739, n_14106, n_14108);
  nand g42291 (n_16337, n_14911, rst_n);
  or g42292 (n_15944, n_15943, wc1193);
  not gc1193 (wc1193, n_14369);
  or g42293 (n_15822, n_15821, wc1194);
  not gc1194 (wc1194, n_13962);
  or g42294 (n_18034, wc1195, n_13816);
  not gc1195 (wc1195, sh_reg_out[28]);
  or g42295 (n_13939, n_16092, wc1196);
  not gc1196 (wc1196, sh_reg_in[5]);
  nand g42296 (n_22075, out_fifo_write_pointer[0], n_14578);
  or g42297 (n_13832, out_fifo_write_pointer[0], n_14578);
  nand g42298 (n_15467, n_22075, n_13832);
  nand g42299 (n_22077, n_14240, n_14277);
  or g42300 (n_22078, n_14240, n_14277);
  nand g42301 (n_14278, n_22077, n_22078);
  or g42302 (n_16124, n_13974, n_13975);
  or g42305 (n_15885, n_15884, wc1197);
  not gc1197 (wc1197, n_14166);
  or g42306 (n_18082, wc1198, n_13816);
  not gc1198 (wc1198, sh_reg_out[17]);
  or g42309 (n_16197, wc1199, n_13924);
  not gc1199 (wc1199, n_13919);
  nand g42312 (n_20811, n_15019, n_14108);
  or g42313 (n_17266, wc1200, n_13816);
  not gc1200 (wc1200, sh_reg_out[16]);
  nand g42314 (n_16196, n_13923, n_14993);
  nand g42315 (n_15777, n_15775, n_15776);
  or g42316 (n_15954, wc1201, n_13944);
  not gc1201 (wc1201, \data_stack_mem[8] [6]);
  nand g42317 (n_14140, n_15656, n_15657);
  nand g42318 (n_15904, n_14275, n_15903);
  nand g42319 (n_15997, n_15502, n_15501);
  or g42320 (n_15926, n_15925, wc1202);
  not gc1202 (wc1202, n_14327);
  nand g42321 (n_15703, n_15490, n_15489);
  or g42322 (n_22082, wc1203, n_14376);
  not gc1203 (wc1203, n_14463);
  or g42323 (n_22083, n_14463, wc1204);
  not gc1204 (wc1204, n_14376);
  nand g42324 (n_14464, n_22082, n_22083);
  nand g42325 (n_16290, n_15509, n_15508);
  nand g42326 (n_15724, n_15515, n_14883);
  or g42327 (n_15966, wc1205, n_13944);
  not gc1205 (wc1205, \data_stack_mem[8] [0]);
  or g42328 (n_14417, wc1206, n_14416);
  not gc1206 (wc1206, n_13875);
  or g42329 (n_13913, sh_reg_in[5], n_13911);
  nand g42330 (n_16043, n_15514, n_15513);
  nand g42331 (n_16006, n_15504, n_15503);
  or g42332 (n_15960, wc1207, n_13944);
  not gc1207 (wc1207, \data_stack_mem[8] [3]);
  or g42333 (n_22084, wc1208, n_14103);
  not gc1208 (wc1208, n_14125);
  or g42334 (n_22085, n_14125, wc1209);
  not gc1209 (wc1209, n_14103);
  nand g42335 (n_14126, n_22084, n_22085);
  or g42336 (n_15821, n_15820, wc1210);
  not gc1210 (wc1210, n_13999);
  nand g42337 (n_16170, n_15507, n_15506);
  or g42338 (n_15799, n_15798, wc1211);
  not gc1211 (wc1211, n_13920);
  nand g42339 (n_15990, n_15498, n_14889);
  nand g42340 (n_15472, n_15686, n_15687);
  or g42341 (n_15951, wc1212, n_13944);
  not gc1212 (wc1212, \data_stack_mem[8] [7]);
  or g42342 (n_14676, sh_reg_in[8], wc1213);
  not gc1213 (wc1213, n_15465);
  nand g42343 (n_15943, n_14461, n_14462);
  nand g42344 (n_15476, n_15695, n_15696);
  or g42345 (n_15788, n_15786, wc1214);
  not gc1214 (wc1214, n_13920);
  nand g42346 (n_22086, out_fifo_read_pointer[0], n_13851);
  or g42347 (n_22087, out_fifo_read_pointer[0], n_13851);
  nand g42348 (n_15484, n_22086, n_22087);
  or g42349 (n_15963, wc1215, n_13944);
  not gc1215 (wc1215, \data_stack_mem[8] [2]);
  or g42350 (n_16089, n_13875, n_13911);
  or g42351 (n_22088, wc1216, n_14307);
  not gc1216 (wc1216, n_14329);
  or g42352 (n_22089, n_14329, wc1217);
  not gc1217 (wc1217, n_14307);
  nand g42353 (n_14330, n_22088, n_22089);
  nand g42354 (n_15985, n_15495, n_15494);
  or g42355 (n_20325, wc1218, n_13910);
  not gc1218 (wc1218, \data_stack_mem[0] [7]);
  or g42356 (n_22090, wc1219, n_14276);
  not gc1219 (wc1219, n_14241);
  or g42357 (n_22091, n_14241, wc1220);
  not gc1220 (wc1220, n_14276);
  nand g42358 (n_14277, n_22090, n_22091);
  or g42359 (n_15863, n_15862, wc1221);
  not gc1221 (wc1221, n_14123);
  or g42360 (n_16092, n_13874, n_13911);
  nand g42361 (n_16165, n_15500, n_15499);
  nand g42362 (n_15765, n_15763, n_15764);
  or g42363 (n_22092, wc1222, n_13973);
  not gc1222 (wc1222, n_14000);
  or g42364 (n_22093, n_14000, wc1223);
  not gc1223 (wc1223, n_13973);
  nand g42365 (n_14001, n_22092, n_22093);
  or g42366 (n_15459, n_15581, n_15582);
  or g42367 (n_13906, n_15017, wc1224);
  not gc1224 (wc1224, rst_n);
  or g42368 (n_15957, wc1225, n_13944);
  not gc1225 (wc1225, \data_stack_mem[8] [4]);
  nand g42369 (n_13816, n_15017, rst_n);
  or g42370 (n_19027, n_15456, sh_reg_in[0]);
  nand g42371 (n_14866, rst_n, n_13853);
  nand g42372 (n_14108, n_15615, n_20808);
  or g42373 (n_22094, wc1226, n_14047);
  not gc1226 (wc1226, n_14024);
  or g42374 (n_22095, n_14024, wc1227);
  not gc1227 (wc1227, n_14047);
  nand g42375 (n_14048, n_22094, n_22095);
  nand g42376 (n_16024, n_14937, n_16023);
  nand g42377 (n_22096, n_15026, n_14173);
  or g42378 (n_22097, n_15026, n_14173);
  nand g42379 (n_14210, n_22096, n_22097);
  or g42380 (n_16086, sh_reg_in[8], wc1228);
  not gc1228 (wc1228, n_15466);
  nand g42381 (n_16032, n_15512, n_15511);
  nand g42382 (n_15975, n_15492, n_15491);
  or g42383 (n_15884, n_15883, wc1229);
  not gc1229 (wc1229, n_14209);
  or g42384 (n_13945, wc1230, n_13944);
  not gc1230 (wc1230, n_13937);
  or g42385 (n_15842, n_15841, wc1231);
  not gc1231 (wc1231, n_14044);
  or g42386 (n_15518, wc1232, n_15729);
  not gc1232 (wc1232, n_13873);
  or g42387 (n_13911, wc1233, n_13871);
  not gc1233 (wc1233, n_13870);
  nand g42388 (n_13923, n_13921, n_15804);
  or g42389 (n_14877, \data_stack_mem[6] [5], n_13916);
  nand g42390 (n_15468, n_14396, n_15678);
  or g42391 (n_14937, n_13916, wc1234);
  not gc1234 (wc1234, \data_stack_mem[6] [0]);
  nand g42392 (n_13910, n_13870, n_13871);
  nand g42393 (n_15502, n_14107, n_15711);
  or g42394 (n_15497, \data_stack_mem[6] [3], n_13916);
  or g42395 (n_16422, \data_stack_mem[0] [7], n_14396);
  or g42396 (n_13944, sh_reg_in[1], n_13943);
  or g42397 (n_14461, n_13916, wc1235);
  not gc1235 (wc1235, \data_stack_mem[6] [7]);
  or g42398 (n_13965, n_13916, wc1236);
  not gc1236 (wc1236, \data_stack_mem[6] [1]);
  or g42399 (n_13851, n_15540, wc1237);
  not gc1237 (wc1237, sh_reg_out_bit_counter[0]);
  nand g42400 (n_14463, n_14380, n_15675);
  or g42401 (n_15763, n_15762, wc1238);
  not gc1238 (wc1238, n_13920);
  nand g42402 (n_15465, n_13855, n_15633);
  or g42403 (n_15764, n_13947, n_13977);
  or g42404 (n_15481, n_13937, wc1239);
  not gc1239 (wc1239, n_15594);
  or g42405 (n_13983, \data_stack_mem[6] [1], n_13916);
  or g42406 (n_15775, n_13922, n_13977);
  or g42407 (n_15776, n_15774, wc1240);
  not gc1240 (wc1240, n_13920);
  nand g42408 (n_15841, n_14046, n_15840);
  nand g42409 (n_14329, n_14311, n_15672);
  nand g42410 (n_14000, n_13977, n_15660);
  or g42411 (n_14327, n_13916, wc1241);
  not gc1241 (wc1241, \data_stack_mem[6] [6]);
  or g42412 (n_14043, n_13940, wc1242);
  not gc1242 (wc1242, n_13937);
  or g42413 (n_14416, wc1243, n_13871);
  not gc1243 (wc1243, n_15651);
  nand g42414 (n_15498, n_15657, n_14029);
  or g42415 (n_15582, n_15579, n_15580);
  nand g42416 (n_15862, n_14124, n_15861);
  or g42417 (n_15787, n_14028, n_14030);
  or g42418 (n_15482, n_13937, wc1244);
  not gc1244 (wc1244, n_15597);
  nand g42419 (n_15786, n_14027, n_14030);
  or g42420 (n_14042, n_13937, n_13940);
  or g42421 (n_14867, wc1245, n_13937);
  not gc1245 (wc1245, sh_reg_in[1]);
  or g42422 (n_14044, n_13916, wc1246);
  not gc1246 (wc1246, \data_stack_mem[6] [2]);
  nand g42423 (n_14047, n_14028, n_15663);
  or g42424 (n_15500, \data_stack_mem[6] [2], n_13916);
  or g42425 (n_15798, n_14064, wc1247);
  not gc1247 (wc1247, n_14027);
  or g42426 (n_15800, n_14028, wc1248);
  not gc1248 (wc1248, n_14064);
  or g42427 (n_15480, n_13937, wc1249);
  not gc1249 (wc1249, n_15591);
  nand g42428 (n_15883, n_14208, n_15882);
  nand g42429 (n_20808, n_15009, n_14030);
  nand g42430 (n_15514, n_14178, n_15717);
  or g42431 (n_14123, n_13916, wc1250);
  not gc1250 (wc1250, \data_stack_mem[6] [3]);
  nand g42432 (n_14125, n_14106, n_15666);
  nand g42433 (n_15466, data_stack_pointer[0], n_14586);
  nand g42434 (n_15656, n_15423, n_14064);
  nand g42435 (n_15512, n_13921, n_13947);
  nand g42436 (n_15686, n_15471, n_15470);
  or g42437 (n_15729, wc1251, n_13871);
  not gc1251 (wc1251, n_13875);
  or g42438 (n_15696, wc1252, n_13828);
  not gc1252 (wc1252, sh_bit_cnt[3]);
  nand g42439 (n_15820, n_13998, n_15819);
  or g42440 (n_14167, \data_stack_mem[6] [4], n_13916);
  nand g42441 (n_14276, n_14244, n_15669);
  or g42442 (n_14166, n_13916, wc1253);
  not gc1253 (wc1253, \data_stack_mem[6] [4]);
  or g42443 (n_14274, n_13916, wc1254);
  not gc1254 (wc1254, \data_stack_mem[6] [5]);
  nand g42444 (n_15026, n_14177, n_14178);
  or g42445 (n_15509, \data_stack_mem[6] [0], n_13916);
  or g42446 (n_15483, n_13937, wc1255);
  not gc1255 (wc1255, n_15600);
  or g42447 (n_15496, \data_stack_mem[6] [7], n_13916);
  nand g42448 (n_15474, n_13815, n_15690);
  nand g42449 (n_15504, n_14381, n_15714);
  nand g42450 (n_15495, n_14312, n_15708);
  or g42451 (n_15493, \data_stack_mem[6] [6], n_13916);
  nand g42452 (n_16110, sh_bit_cnt[3], n_13828);
  or g42453 (n_15475, n_13937, wc1256);
  not gc1256 (wc1256, n_15585);
  nand g42454 (n_15469, n_14396, n_15681);
  or g42455 (n_16428, wc1257, n_14396);
  not gc1257 (wc1257, \data_stack_mem[0] [7]);
  nand g42456 (n_15925, n_14328, n_15924);
  nand g42457 (n_16232, sh_reg_out_bit_counter[4], n_13815);
  nand g42458 (n_15924, \data_stack_mem[1] [6], n_13920);
  or g42459 (n_20170, wc1258, n_13873);
  not gc1258 (wc1258, \data_stack_mem[0] [6]);
  nand g42460 (n_13916, n_13914, n_15450);
  nand g42461 (n_15681, \data_stack_mem[0] [7], n_13920);
  nand g42462 (n_14396, n_13920, \data_stack_mem[1] [7]);
  or g42463 (n_14029, wc1259, n_13920);
  not gc1259 (wc1259, \data_stack_mem[0] [2]);
  or g42464 (n_15494, \data_stack_mem[5] [6], n_13917);
  nand g42465 (n_15690, sh_reg_out_bit_counter[3], n_13814);
  or g42466 (n_20290, wc1260, n_13873);
  not gc1260 (wc1260, \data_stack_mem[0] [7]);
  nand g42467 (n_15473, n_13814, n_15639);
  or g42468 (n_15651, sh_reg_in[5], wc1261);
  not gc1261 (wc1261, n_13940);
  or g42469 (n_14252, \data_stack_mem[5] [5], n_13917);
  or g42470 (n_19155, wc1262, n_13873);
  not gc1262 (wc1262, \data_stack_mem[0] [0]);
  nand g42471 (n_15580, n_15575, n_15576);
  nand g42472 (n_16467, n_15457, rst_n);
  nand g42473 (n_16023, n_15505, n_13920);
  or g42474 (n_14244, wc1263, n_14243);
  not gc1263 (wc1263, n_13920);
  or g42475 (n_13921, wc1264, n_13920);
  not gc1264 (wc1264, \data_stack_mem[0] [0]);
  nand g42476 (n_13918, n_13914, n_15630);
  or g42477 (n_14872, wc1265, n_13920);
  not gc1265 (wc1265, \data_stack_mem[0] [5]);
  or g42478 (n_14236, n_13917, wc1266);
  not gc1266 (wc1266, \data_stack_mem[5] [5]);
  or g42479 (n_15660, \data_stack_mem[0] [1], n_13920);
  or g42480 (n_14328, n_13917, wc1267);
  not gc1267 (wc1267, \data_stack_mem[5] [6]);
  or g42481 (n_13998, n_13917, wc1268);
  not gc1268 (wc1268, \data_stack_mem[5] [1]);
  or g42482 (n_15672, \data_stack_mem[0] [6], n_13920);
  or g42483 (n_14380, wc1269, n_14378);
  not gc1269 (wc1269, n_13920);
  or g42484 (n_14209, n_13917, wc1270);
  not gc1270 (wc1270, \data_stack_mem[5] [4]);
  nand g42485 (n_13875, n_13874, sh_reg_in[5]);
  or g42486 (n_15506, \data_stack_mem[5] [0], n_13917);
  or g42487 (n_13850, n_15528, wc1271);
  not gc1271 (wc1271, rst_n);
  nand g42488 (n_15774, n_13976, n_13922);
  or g42489 (n_13871, sh_reg_in[6], n_15546);
  nand g42490 (n_15579, n_15573, n_15574);
  nand g42491 (n_15840, \data_stack_mem[1] [2], n_13920);
  or g42492 (n_15669, \data_stack_mem[0] [5], n_13920);
  nand g42493 (n_15819, \data_stack_mem[1] [1], n_13920);
  or g42494 (n_15501, \data_stack_mem[5] [3], n_13917);
  or g42495 (n_15678, \data_stack_mem[0] [7], wc1272);
  not gc1272 (wc1272, n_13920);
  nand g42496 (n_14177, n_14176, n_13920);
  nand g42497 (n_15581, n_15577, n_15578);
  or g42498 (n_19564, wc1273, n_13873);
  not gc1273 (wc1273, \data_stack_mem[0] [2]);
  nand g42499 (n_15695, sh_bit_cnt[2], n_14912);
  nand g42500 (n_15903, \data_stack_mem[1] [5], n_13920);
  nand g42501 (n_15471, n_14912, n_15636);
  or g42502 (n_14879, \data_stack_mem[5] [4], n_13917);
  or g42503 (n_14586, data_stack_pointer[1], wc1274);
  not gc1274 (wc1274, n_15519);
  or g42504 (n_15666, \data_stack_mem[0] [3], n_13920);
  or g42505 (n_14124, n_13917, wc1275);
  not gc1275 (wc1275, \data_stack_mem[5] [3]);
  or g42506 (n_13977, wc1276, n_13976);
  not gc1276 (wc1276, n_13920);
  or g42507 (n_14951, n_13917, wc1277);
  not gc1277 (wc1277, \data_stack_mem[5] [0]);
  or g42508 (n_14388, \data_stack_mem[5] [7], n_13917);
  or g42509 (n_14106, wc1278, n_14105);
  not gc1278 (wc1278, n_13920);
  nand g42510 (n_15762, n_13947, n_13976);
  or g42511 (n_14107, wc1279, n_13920);
  not gc1279 (wc1279, \data_stack_mem[0] [3]);
  or g42512 (n_14312, wc1280, n_13920);
  not gc1280 (wc1280, \data_stack_mem[0] [6]);
  nand g42513 (n_15882, \data_stack_mem[1] [4], n_13920);
  or g42514 (n_19942, wc1281, n_13873);
  not gc1281 (wc1281, \data_stack_mem[0] [4]);
  or g42515 (n_14311, wc1282, n_14310);
  not gc1282 (wc1282, n_13920);
  or g42516 (n_14871, wc1283, n_13920);
  not gc1283 (wc1283, \data_stack_mem[0] [1]);
  nand g42517 (n_14064, n_15611, n_15612);
  nand g42518 (n_15633, n_15464, rst_n);
  or g42519 (n_15499, \data_stack_mem[5] [2], n_13917);
  or g42520 (n_15663, \data_stack_mem[0] [2], n_13920);
  or g42521 (n_14045, n_13917, wc1284);
  not gc1284 (wc1284, \data_stack_mem[5] [2]);
  or g42522 (n_14369, n_13917, wc1285);
  not gc1285 (wc1285, \data_stack_mem[5] [7]);
  or g42523 (n_15492, \data_stack_mem[5] [1], n_13917);
  nand g42524 (n_15804, n_15305, n_13920);
  or g42525 (n_19717, wc1286, n_13873);
  not gc1286 (wc1286, \data_stack_mem[0] [3]);
  or g42526 (n_15675, \data_stack_mem[0] [7], n_13920);
  or g42527 (n_15540, sh_reg_out_bit_counter[4], n_15539);
  nand g42528 (n_13943, n_15517, sh_reg_in[0]);
  nand g42529 (n_14030, n_15605, n_15606);
  or g42530 (n_14381, wc1287, n_13920);
  not gc1287 (wc1287, \data_stack_mem[0] [7]);
  or g42531 (n_14028, wc1288, n_14027);
  not gc1288 (wc1288, n_13920);
  nand g42532 (n_13937, data_stack_pointer[3], n_20802);
  nand g42533 (n_15861, \data_stack_mem[1] [3], n_13920);
  or g42534 (n_15630, data_stack_pointer[1], n_13868);
  nand g42535 (n_20256, n_13872, \data_stack_mem[0] [7]);
  or g42536 (n_16452, n_13855, wc1289);
  not gc1289 (wc1289, n_14607);
  nand g42537 (n_14240, \data_stack_mem[3] [5], n_13914);
  or g42538 (n_14239, wc1290, \data_stack_mem[3] [5]);
  not gc1290 (wc1290, n_13914);
  nand g42539 (n_14243, n_14995, n_15624);
  nand g42540 (n_13873, n_13872, sh_reg_in[4]);
  nand g42541 (n_15639, sh_reg_out_bit_counter[2], n_13813);
  nand g42542 (n_13917, n_13914, n_15446);
  nand g42543 (n_15457, n_14607, n_15552);
  or g42544 (n_15546, sh_reg_in[3], n_15545);
  or g42545 (n_20835, n_13855, wc1291);
  not gc1291 (wc1291, n_13868);
  nand g42546 (n_15528, n_15526, n_15527);
  or g42547 (n_15450, data_stack_pointer[3], wc1292);
  not gc1292 (wc1292, n_13915);
  nand g42548 (n_14172, \data_stack_mem[3] [4], n_13914);
  or g42549 (n_14171, wc1293, \data_stack_mem[3] [4]);
  not gc1293 (wc1293, n_13914);
  nand g42550 (n_14176, n_15041, n_15621);
  nand g42551 (n_15477, n_13813, n_15588);
  or g42552 (n_15510, \data_stack_mem[3] [0], wc1294);
  not gc1294 (wc1294, n_13914);
  or g42553 (n_15519, data_stack_pointer[2], n_14585);
  nand g42554 (n_14102, \data_stack_mem[3] [3], n_13914);
  or g42555 (n_14101, wc1295, \data_stack_mem[3] [3]);
  not gc1295 (wc1295, n_13914);
  nand g42556 (n_14105, n_15019, n_15618);
  nand g42557 (n_14310, n_14989, n_15627);
  or g42558 (n_14987, wc1296, n_13914);
  not gc1296 (wc1296, data_stack_pointer[0]);
  or g42559 (n_15611, wc1297, n_13947);
  not gc1297 (wc1297, n_15415);
  or g42560 (n_14305, wc1298, \data_stack_mem[3] [6]);
  not gc1298 (wc1298, n_13914);
  nand g42561 (n_14046, \data_stack_mem[3] [2], n_13914);
  or g42562 (n_14889, wc1299, \data_stack_mem[3] [2]);
  not gc1299 (wc1299, n_13914);
  or g42563 (n_14372, wc1300, \data_stack_mem[3] [7]);
  not gc1300 (wc1300, n_13914);
  nand g42564 (n_14306, \data_stack_mem[3] [6], n_13914);
  nand g42565 (n_15605, n_13922, n_14975);
  nand g42566 (n_14027, n_15009, n_15615);
  or g42567 (n_15576, n_13825, wc1301);
  not gc1301 (wc1301, n_13902);
  or g42568 (n_15575, wc1302, n_14909);
  not gc1302 (wc1302, n_13904);
  nand g42569 (n_14373, \data_stack_mem[3] [7], n_13914);
  or g42570 (n_15574, wc1303, n_15038);
  not gc1303 (wc1303, n_13903);
  nand g42571 (n_13972, \data_stack_mem[3] [1], n_13914);
  or g42572 (n_13971, wc1304, \data_stack_mem[3] [1]);
  not gc1304 (wc1304, n_13914);
  or g42573 (n_15577, n_13839, wc1305);
  not gc1305 (wc1305, n_13905);
  nand g42574 (n_13976, n_14975, n_15606);
  or g42575 (n_15464, data_stack_pointer[1], n_14585);
  or g42576 (n_15539, sh_reg_out_bit_counter[3], n_15538);
  nand g42577 (n_15517, data_stack_pointer[3], n_15531);
  or g42578 (n_20802, data_stack_pointer[0], n_15531);
  or g42579 (n_13919, n_13914, wc1306);
  not gc1306 (wc1306, n_13915);
  nand g42580 (n_15305, n_13922, n_15549);
  or g42581 (n_13920, data_stack_pointer[1], n_13914);
  nand g42582 (n_14980, \data_stack_mem[3] [0], n_13914);
  or g42583 (n_16317, data_stack_pointer[2], wc1307);
  not gc1307 (wc1307, n_14585);
  nand g42584 (n_13915, data_stack_pointer[0], data_stack_pointer[1]);
  or g42585 (n_13914, data_stack_pointer[2], data_stack_pointer[3]);
  or g42586 (n_15549, wc1308, \data_stack_mem[1] [0]);
  not gc1308 (wc1308, \data_stack_mem[0] [0]);
  or g42587 (n_13905, wc1309, out_fifo_read_pointer[2]);
  not gc1309 (wc1309, out_fifo_read_pointer[1]);
  or g42588 (n_13904, out_fifo_read_pointer[1], wc1310);
  not gc1310 (wc1310, out_fifo_read_pointer[2]);
  or g42589 (n_13903, out_fifo_read_pointer[2],
       out_fifo_read_pointer[1]);
  nand g42590 (n_13902, out_fifo_read_pointer[2],
       out_fifo_read_pointer[1]);
  or g42591 (n_13942, wc1311, sh_reg_in[4]);
  not gc1311 (wc1311, sh_reg_in[1]);
  or g42592 (n_15531, data_stack_pointer[1], data_stack_pointer[2]);
  nand g42593 (n_13947, \data_stack_mem[0] [0], \data_stack_mem[1] [0]);
  or g42594 (n_15606, wc1312, \data_stack_mem[1] [1]);
  not gc1312 (wc1312, \data_stack_mem[0] [1]);
  or g42595 (n_15615, wc1313, \data_stack_mem[1] [2]);
  not gc1313 (wc1313, \data_stack_mem[0] [2]);
  nand g42596 (n_15612, \data_stack_mem[0] [1], \data_stack_mem[1] [1]);
  or g42597 (n_15618, wc1314, \data_stack_mem[1] [3]);
  not gc1314 (wc1314, \data_stack_mem[0] [3]);
  nand g42598 (n_15657, \data_stack_mem[0] [2], \data_stack_mem[1] [2]);
  or g42599 (n_15621, wc1315, \data_stack_mem[1] [4]);
  not gc1315 (wc1315, \data_stack_mem[0] [4]);
  nand g42600 (n_15711, \data_stack_mem[0] [3], \data_stack_mem[1] [3]);
  or g42601 (n_15545, sh_reg_in[2], sh_reg_in[7]);
  or g42602 (n_15624, wc1316, \data_stack_mem[1] [5]);
  not gc1316 (wc1316, \data_stack_mem[0] [5]);
  nand g42603 (n_15717, \data_stack_mem[0] [4], \data_stack_mem[1] [4]);
  nand g42604 (n_13855, rst_n, data_stack_pointer[2]);
  or g42605 (n_15627, wc1317, \data_stack_mem[1] [6]);
  not gc1317 (wc1317, \data_stack_mem[0] [6]);
  nand g42606 (n_16191, \data_stack_mem[0] [5], \data_stack_mem[1] [5]);
  or g42607 (n_22098, wc1318, \data_stack_mem[1] [7]);
  not gc1318 (wc1318, \data_stack_mem[0] [7]);
  or g42608 (n_22099, \data_stack_mem[0] [7], wc1319);
  not gc1319 (wc1319, \data_stack_mem[1] [7]);
  nand g42609 (n_14378, n_22098, n_22099);
  nand g42610 (n_15708, \data_stack_mem[0] [6], \data_stack_mem[1] [6]);
  or g42611 (n_15594, \data_stack_mem[8] [2], wc1320);
  not gc1320 (wc1320, sh_reg_in[0]);
  or g42612 (n_15591, \data_stack_mem[8] [4], wc1321);
  not gc1321 (wc1321, sh_reg_in[0]);
  nand g42613 (n_20301, \data_stack_mem[0] [7], sh_reg_in[4]);
  or g42614 (n_15600, \data_stack_mem[8] [7], wc1322);
  not gc1322 (wc1322, sh_reg_in[0]);
  nand g42615 (n_15714, \data_stack_mem[0] [7], \data_stack_mem[1] [7]);
  or g42616 (n_15585, \data_stack_mem[8] [6], wc1323);
  not gc1323 (wc1323, sh_reg_in[0]);
  or g42617 (n_15597, \data_stack_mem[8] [3], wc1324);
  not gc1324 (wc1324, sh_reg_in[0]);
  nand g42618 (n_14585, data_stack_pointer[0], data_stack_pointer[3]);
  or g42619 (n_15538, sh_reg_out_bit_counter[1],
       sh_reg_out_bit_counter[2]);
  or g42620 (n_15578, wc1325, out_fifo_write_pointer[0]);
  not gc1325 (wc1325, out_fifo_read_pointer[0]);
  or g42621 (n_15573, out_fifo_read_pointer[0], wc1326);
  not gc1326 (wc1326, out_fifo_write_pointer[0]);
  nand g42622 (n_15636, sh_bit_cnt[0], sh_bit_cnt[1]);
  nand g42623 (n_15687, sh_bit_cnt[1], enable_n);
  nand g42624 (n_15588, sh_reg_out_bit_counter[0],
       sh_reg_out_bit_counter[1]);
  or g42625 (n_15526, sh_bit_cnt[0], enable_n);
  nand g42626 (n_15527, sh_bit_cnt[0], enable_n);
  or g42627 (n_15552, data_stack_pointer[0], wc1327);
  not gc1327 (wc1327, data_stack_pointer[3]);
  or g42628 (n_16443, data_stack_pointer[3], wc1328);
  not gc1328 (wc1328, rst_n);
  or g42629 (n_16458, data_stack_pointer[0], wc1329);
  not gc1329 (wc1329, rst_n);
  and g42630 (n_22052, n_15476, rst_n);
  and g42631 (n_22053, wc1330, sh_reg_out[22]);
  not gc1330 (wc1330, n_13816);
  and g42632 (n_22054, n_15477, wc1331);
  not gc1331 (wc1331, n_13816);
  and g42633 (n_22060, wc1332, sh_reg_out[21]);
  not gc1332 (wc1332, n_13816);
  and g42634 (n_22061, wc1333, sh_reg_out[18]);
  not gc1333 (wc1333, n_13816);
  and g42635 (n_22062, wc1334, sh_reg_out[25]);
  not gc1334 (wc1334, n_13816);
  and g42636 (n_22073, wc1335, sh_reg_out[8]);
  not gc1335 (wc1335, n_13816);
  and g42637 (n_22074, wc1336, sh_reg_out[26]);
  not gc1336 (wc1336, n_13816);
  and g42638 (n_22079, wc1337, sh_reg_out[24]);
  not gc1337 (wc1337, n_13816);
  and g42639 (n_22080, wc1338, sh_reg_out[23]);
  not gc1338 (wc1338, n_13816);
  and g42640 (n_22081, n_15472, rst_n);
  and g42641 (n_22055, n_15484, rst_n);
  and g42642 (n_22038, n_15485, rst_n);
  and g42643 (n_22039, n_15467, rst_n);
  and g42644 (n_22018, n_15486, rst_n);
  and g42645 (n_22029, n_15461, rst_n);
  and g42646 (n_22001, n_15460, rst_n);
  or g42650 (n_14525, wc1339, n_14524);
  not gc1339 (wc1339, n_15030);
  or g42651 (n_14526, wc1340, n_14525);
  not gc1340 (wc1340, n_14998);
  CDN_flop \out_fifo_read_pointer_reg[0] (.clk (clk), .d (n_22055),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[0]));
  CDN_flop \out_fifo_read_pointer_reg[1] (.clk (clk), .d (n_22038),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[1]));
  CDN_flop \out_fifo_read_pointer_reg[2] (.clk (clk), .d (n_22018),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[2]));
  CDN_flop \out_fifo_reg[0][0][0] (.clk (clk), .d (n_14559), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [0]));
  CDN_flop \out_fifo_reg[0][0][1] (.clk (clk), .d (n_13959), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [1]));
  CDN_flop \out_fifo_reg[0][0][2] (.clk (clk), .d (n_14090), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [2]));
  CDN_flop \out_fifo_reg[0][0][3] (.clk (clk), .d (n_14091), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [3]));
  CDN_flop \out_fifo_reg[0][0][4] (.clk (clk), .d (n_14162), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [4]));
  CDN_flop \out_fifo_reg[0][0][5] (.clk (clk), .d (n_14230), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [5]));
  CDN_flop \out_fifo_reg[0][0][6] (.clk (clk), .d (n_14296), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [6]));
  CDN_flop \out_fifo_reg[0][0][7] (.clk (clk), .d (n_14365), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [7]));
  CDN_flop \out_fifo_reg[0][0][8] (.clk (clk), .d (n_14489), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [8]));
  CDN_flop \out_fifo_reg[0][1][0] (.clk (clk), .d (n_14670), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [0]));
  CDN_flop \out_fifo_reg[0][1][1] (.clk (clk), .d (n_14488), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [1]));
  CDN_flop \out_fifo_reg[0][1][2] (.clk (clk), .d (n_14520), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [2]));
  CDN_flop \out_fifo_reg[0][1][3] (.clk (clk), .d (n_14558), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [3]));
  CDN_flop \out_fifo_reg[0][1][4] (.clk (clk), .d (n_14534), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [4]));
  CDN_flop \out_fifo_reg[0][1][5] (.clk (clk), .d (n_14708), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [5]));
  CDN_flop \out_fifo_reg[0][1][6] (.clk (clk), .d (n_14707), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [6]));
  CDN_flop \out_fifo_reg[0][1][7] (.clk (clk), .d (n_14709), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [7]));
  CDN_flop \out_fifo_reg[0][1][8] (.clk (clk), .d (n_14706), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [8]));
  CDN_flop \out_fifo_reg[0][2][0] (.clk (clk), .d (n_13898), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [0]));
  CDN_flop \out_fifo_reg[0][2][1] (.clk (clk), .d (n_14574), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [1]));
  CDN_flop \out_fifo_reg[0][2][8] (.clk (clk), .d (n_14575), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [8]));
  CDN_flop \out_fifo_reg[0][2][9] (.clk (clk), .d (1'b1), .sena
       (n_13847), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (\out_fifo[0][2] [9]));
  CDN_flop \out_fifo_reg[1][0][0] (.clk (clk), .d (n_14551), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [0]));
  CDN_flop \out_fifo_reg[1][0][1] (.clk (clk), .d (n_13955), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [1]));
  CDN_flop \out_fifo_reg[1][0][2] (.clk (clk), .d (n_14082), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [2]));
  CDN_flop \out_fifo_reg[1][0][3] (.clk (clk), .d (n_14083), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [3]));
  CDN_flop \out_fifo_reg[1][0][4] (.clk (clk), .d (n_14158), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [4]));
  CDN_flop \out_fifo_reg[1][0][5] (.clk (clk), .d (n_14226), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [5]));
  CDN_flop \out_fifo_reg[1][0][6] (.clk (clk), .d (n_14292), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [6]));
  CDN_flop \out_fifo_reg[1][0][7] (.clk (clk), .d (n_14361), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [7]));
  CDN_flop \out_fifo_reg[1][0][8] (.clk (clk), .d (n_14481), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [8]));
  CDN_flop \out_fifo_reg[1][1][0] (.clk (clk), .d (n_14666), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [0]));
  CDN_flop \out_fifo_reg[1][1][1] (.clk (clk), .d (n_14480), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [1]));
  CDN_flop \out_fifo_reg[1][1][2] (.clk (clk), .d (n_14516), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [2]));
  CDN_flop \out_fifo_reg[1][1][3] (.clk (clk), .d (n_14550), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [3]));
  CDN_flop \out_fifo_reg[1][1][4] (.clk (clk), .d (n_14530), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [4]));
  CDN_flop \out_fifo_reg[1][1][5] (.clk (clk), .d (n_14734), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [5]));
  CDN_flop \out_fifo_reg[1][1][6] (.clk (clk), .d (n_14733), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [6]));
  CDN_flop \out_fifo_reg[1][1][7] (.clk (clk), .d (n_14731), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [7]));
  CDN_flop \out_fifo_reg[1][1][8] (.clk (clk), .d (n_14732), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [8]));
  CDN_flop \out_fifo_reg[1][2][0] (.clk (clk), .d (n_13886), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [0]));
  CDN_flop \out_fifo_reg[1][2][1] (.clk (clk), .d (n_14566), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [1]));
  CDN_flop \out_fifo_reg[1][2][8] (.clk (clk), .d (n_14567), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [8]));
  CDN_flop \out_fifo_reg[1][2][9] (.clk (clk), .d (1'b1), .sena
       (n_13845), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (\out_fifo[1][2] [9]));
  CDN_flop \out_fifo_reg[2][0][0] (.clk (clk), .d (n_14549), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [0]));
  CDN_flop \out_fifo_reg[2][0][1] (.clk (clk), .d (n_13954), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [1]));
  CDN_flop \out_fifo_reg[2][0][2] (.clk (clk), .d (n_14080), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [2]));
  CDN_flop \out_fifo_reg[2][0][3] (.clk (clk), .d (n_14081), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [3]));
  CDN_flop \out_fifo_reg[2][0][4] (.clk (clk), .d (n_14157), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [4]));
  CDN_flop \out_fifo_reg[2][0][5] (.clk (clk), .d (n_14225), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [5]));
  CDN_flop \out_fifo_reg[2][0][6] (.clk (clk), .d (n_14291), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [6]));
  CDN_flop \out_fifo_reg[2][0][7] (.clk (clk), .d (n_14360), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [7]));
  CDN_flop \out_fifo_reg[2][0][8] (.clk (clk), .d (n_14479), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [8]));
  CDN_flop \out_fifo_reg[2][1][0] (.clk (clk), .d (n_14665), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [0]));
  CDN_flop \out_fifo_reg[2][1][1] (.clk (clk), .d (n_14478), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [1]));
  CDN_flop \out_fifo_reg[2][1][2] (.clk (clk), .d (n_14515), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [2]));
  CDN_flop \out_fifo_reg[2][1][3] (.clk (clk), .d (n_14548), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [3]));
  CDN_flop \out_fifo_reg[2][1][4] (.clk (clk), .d (n_14529), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [4]));
  CDN_flop \out_fifo_reg[2][1][5] (.clk (clk), .d (n_14724), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [5]));
  CDN_flop \out_fifo_reg[2][1][6] (.clk (clk), .d (n_14723), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [6]));
  CDN_flop \out_fifo_reg[2][1][7] (.clk (clk), .d (n_14722), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [7]));
  CDN_flop \out_fifo_reg[2][1][8] (.clk (clk), .d (n_14721), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [8]));
  CDN_flop \out_fifo_reg[2][2][0] (.clk (clk), .d (n_13883), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [0]));
  CDN_flop \out_fifo_reg[2][2][1] (.clk (clk), .d (n_14564), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [1]));
  CDN_flop \out_fifo_reg[2][2][8] (.clk (clk), .d (n_14565), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [8]));
  CDN_flop \out_fifo_reg[2][2][9] (.clk (clk), .d (1'b1), .sena
       (n_13843), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (\out_fifo[2][2] [9]));
  CDN_flop \out_fifo_reg[3][0][0] (.clk (clk), .d (n_14555), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [0]));
  CDN_flop \out_fifo_reg[3][0][1] (.clk (clk), .d (n_13957), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [1]));
  CDN_flop \out_fifo_reg[3][0][2] (.clk (clk), .d (n_14086), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [2]));
  CDN_flop \out_fifo_reg[3][0][3] (.clk (clk), .d (n_14087), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [3]));
  CDN_flop \out_fifo_reg[3][0][4] (.clk (clk), .d (n_14160), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [4]));
  CDN_flop \out_fifo_reg[3][0][5] (.clk (clk), .d (n_14228), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [5]));
  CDN_flop \out_fifo_reg[3][0][6] (.clk (clk), .d (n_14294), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [6]));
  CDN_flop \out_fifo_reg[3][0][7] (.clk (clk), .d (n_14363), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [7]));
  CDN_flop \out_fifo_reg[3][0][8] (.clk (clk), .d (n_14485), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [8]));
  CDN_flop \out_fifo_reg[3][1][0] (.clk (clk), .d (n_14668), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [0]));
  CDN_flop \out_fifo_reg[3][1][1] (.clk (clk), .d (n_14484), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [1]));
  CDN_flop \out_fifo_reg[3][1][2] (.clk (clk), .d (n_14518), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [2]));
  CDN_flop \out_fifo_reg[3][1][3] (.clk (clk), .d (n_14554), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [3]));
  CDN_flop \out_fifo_reg[3][1][4] (.clk (clk), .d (n_14532), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [4]));
  CDN_flop \out_fifo_reg[3][1][5] (.clk (clk), .d (n_14741), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [5]));
  CDN_flop \out_fifo_reg[3][1][6] (.clk (clk), .d (n_14743), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [6]));
  CDN_flop \out_fifo_reg[3][1][7] (.clk (clk), .d (n_14742), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [7]));
  CDN_flop \out_fifo_reg[3][1][8] (.clk (clk), .d (n_14744), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [8]));
  CDN_flop \out_fifo_reg[3][2][0] (.clk (clk), .d (n_13892), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [0]));
  CDN_flop \out_fifo_reg[3][2][1] (.clk (clk), .d (n_14570), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [1]));
  CDN_flop \out_fifo_reg[3][2][8] (.clk (clk), .d (n_14571), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [8]));
  CDN_flop \out_fifo_reg[3][2][9] (.clk (clk), .d (1'b1), .sena
       (n_13841), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (\out_fifo[3][2] [9]));
  CDN_flop \out_fifo_reg[4][0][0] (.clk (clk), .d (n_14561), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [0]));
  CDN_flop \out_fifo_reg[4][0][1] (.clk (clk), .d (n_13960), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [1]));
  CDN_flop \out_fifo_reg[4][0][2] (.clk (clk), .d (n_14092), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [2]));
  CDN_flop \out_fifo_reg[4][0][3] (.clk (clk), .d (n_14093), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [3]));
  CDN_flop \out_fifo_reg[4][0][4] (.clk (clk), .d (n_14163), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [4]));
  CDN_flop \out_fifo_reg[4][0][5] (.clk (clk), .d (n_14231), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [5]));
  CDN_flop \out_fifo_reg[4][0][6] (.clk (clk), .d (n_14297), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [6]));
  CDN_flop \out_fifo_reg[4][0][7] (.clk (clk), .d (n_14366), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [7]));
  CDN_flop \out_fifo_reg[4][0][8] (.clk (clk), .d (n_14491), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [8]));
  CDN_flop \out_fifo_reg[4][1][0] (.clk (clk), .d (n_14671), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [0]));
  CDN_flop \out_fifo_reg[4][1][1] (.clk (clk), .d (n_14490), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [1]));
  CDN_flop \out_fifo_reg[4][1][2] (.clk (clk), .d (n_14521), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [2]));
  CDN_flop \out_fifo_reg[4][1][3] (.clk (clk), .d (n_14560), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [3]));
  CDN_flop \out_fifo_reg[4][1][4] (.clk (clk), .d (n_14535), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [4]));
  CDN_flop \out_fifo_reg[4][1][5] (.clk (clk), .d (n_14716), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [5]));
  CDN_flop \out_fifo_reg[4][1][6] (.clk (clk), .d (n_14717), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [6]));
  CDN_flop \out_fifo_reg[4][1][7] (.clk (clk), .d (n_14719), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [7]));
  CDN_flop \out_fifo_reg[4][1][8] (.clk (clk), .d (n_14718), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [8]));
  CDN_flop \out_fifo_reg[4][2][0] (.clk (clk), .d (n_13901), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [0]));
  CDN_flop \out_fifo_reg[4][2][1] (.clk (clk), .d (n_14576), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [1]));
  CDN_flop \out_fifo_reg[4][2][8] (.clk (clk), .d (n_14577), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [8]));
  CDN_flop \out_fifo_reg[4][2][9] (.clk (clk), .d (1'b1), .sena
       (n_13838), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (\out_fifo[4][2] [9]));
  CDN_flop \out_fifo_reg[5][0][0] (.clk (clk), .d (n_14547), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [0]));
  CDN_flop \out_fifo_reg[5][0][1] (.clk (clk), .d (n_13953), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [1]));
  CDN_flop \out_fifo_reg[5][0][2] (.clk (clk), .d (n_14014), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [2]));
  CDN_flop \out_fifo_reg[5][0][3] (.clk (clk), .d (n_14079), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [3]));
  CDN_flop \out_fifo_reg[5][0][4] (.clk (clk), .d (n_14156), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [4]));
  CDN_flop \out_fifo_reg[5][0][5] (.clk (clk), .d (n_14224), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [5]));
  CDN_flop \out_fifo_reg[5][0][6] (.clk (clk), .d (n_14290), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [6]));
  CDN_flop \out_fifo_reg[5][0][7] (.clk (clk), .d (n_14359), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [7]));
  CDN_flop \out_fifo_reg[5][0][8] (.clk (clk), .d (n_14477), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [8]));
  CDN_flop \out_fifo_reg[5][1][0] (.clk (clk), .d (n_14664), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [0]));
  CDN_flop \out_fifo_reg[5][1][1] (.clk (clk), .d (n_14459), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [1]));
  CDN_flop \out_fifo_reg[5][1][2] (.clk (clk), .d (n_14514), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [2]));
  CDN_flop \out_fifo_reg[5][1][3] (.clk (clk), .d (n_14540), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [3]));
  CDN_flop \out_fifo_reg[5][1][4] (.clk (clk), .d (n_14528), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [4]));
  CDN_flop \out_fifo_reg[5][1][5] (.clk (clk), .d (n_14713), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [5]));
  CDN_flop \out_fifo_reg[5][1][6] (.clk (clk), .d (n_14712), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [6]));
  CDN_flop \out_fifo_reg[5][1][7] (.clk (clk), .d (n_14714), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [7]));
  CDN_flop \out_fifo_reg[5][1][8] (.clk (clk), .d (n_14711), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [8]));
  CDN_flop \out_fifo_reg[5][2][0] (.clk (clk), .d (n_13880), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [0]));
  CDN_flop \out_fifo_reg[5][2][1] (.clk (clk), .d (n_14562), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [1]));
  CDN_flop \out_fifo_reg[5][2][8] (.clk (clk), .d (n_14563), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [8]));
  CDN_flop \out_fifo_reg[5][2][9] (.clk (clk), .d (1'b1), .sena
       (n_13836), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (\out_fifo[5][2] [9]));
  CDN_flop \out_fifo_reg[6][0][0] (.clk (clk), .d (n_14553), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [0]));
  CDN_flop \out_fifo_reg[6][0][1] (.clk (clk), .d (n_13956), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [1]));
  CDN_flop \out_fifo_reg[6][0][2] (.clk (clk), .d (n_14084), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [2]));
  CDN_flop \out_fifo_reg[6][0][3] (.clk (clk), .d (n_14085), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [3]));
  CDN_flop \out_fifo_reg[6][0][4] (.clk (clk), .d (n_14159), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [4]));
  CDN_flop \out_fifo_reg[6][0][5] (.clk (clk), .d (n_14227), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [5]));
  CDN_flop \out_fifo_reg[6][0][6] (.clk (clk), .d (n_14293), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [6]));
  CDN_flop \out_fifo_reg[6][0][7] (.clk (clk), .d (n_14362), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [7]));
  CDN_flop \out_fifo_reg[6][0][8] (.clk (clk), .d (n_14483), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [8]));
  CDN_flop \out_fifo_reg[6][1][0] (.clk (clk), .d (n_14667), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [0]));
  CDN_flop \out_fifo_reg[6][1][1] (.clk (clk), .d (n_14482), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [1]));
  CDN_flop \out_fifo_reg[6][1][2] (.clk (clk), .d (n_14517), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [2]));
  CDN_flop \out_fifo_reg[6][1][3] (.clk (clk), .d (n_14552), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [3]));
  CDN_flop \out_fifo_reg[6][1][4] (.clk (clk), .d (n_14531), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [4]));
  CDN_flop \out_fifo_reg[6][1][5] (.clk (clk), .d (n_14738), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [5]));
  CDN_flop \out_fifo_reg[6][1][6] (.clk (clk), .d (n_14736), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [6]));
  CDN_flop \out_fifo_reg[6][1][7] (.clk (clk), .d (n_14737), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [7]));
  CDN_flop \out_fifo_reg[6][1][8] (.clk (clk), .d (n_14739), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [8]));
  CDN_flop \out_fifo_reg[6][2][0] (.clk (clk), .d (n_13889), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [0]));
  CDN_flop \out_fifo_reg[6][2][1] (.clk (clk), .d (n_14568), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [1]));
  CDN_flop \out_fifo_reg[6][2][8] (.clk (clk), .d (n_14569), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [8]));
  CDN_flop \out_fifo_reg[6][2][9] (.clk (clk), .d (1'b1), .sena
       (n_13834), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (\out_fifo[6][2] [9]));
  CDN_flop \out_fifo_reg[7][0][0] (.clk (clk), .d (n_14557), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [0]));
  CDN_flop \out_fifo_reg[7][0][1] (.clk (clk), .d (n_13958), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [1]));
  CDN_flop \out_fifo_reg[7][0][2] (.clk (clk), .d (n_14088), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [2]));
  CDN_flop \out_fifo_reg[7][0][3] (.clk (clk), .d (n_14089), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [3]));
  CDN_flop \out_fifo_reg[7][0][4] (.clk (clk), .d (n_14161), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [4]));
  CDN_flop \out_fifo_reg[7][0][5] (.clk (clk), .d (n_14229), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [5]));
  CDN_flop \out_fifo_reg[7][0][6] (.clk (clk), .d (n_14295), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [6]));
  CDN_flop \out_fifo_reg[7][0][7] (.clk (clk), .d (n_14364), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [7]));
  CDN_flop \out_fifo_reg[7][0][8] (.clk (clk), .d (n_14487), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [8]));
  CDN_flop \out_fifo_reg[7][1][0] (.clk (clk), .d (n_14669), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [0]));
  CDN_flop \out_fifo_reg[7][1][1] (.clk (clk), .d (n_14486), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [1]));
  CDN_flop \out_fifo_reg[7][1][2] (.clk (clk), .d (n_14519), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [2]));
  CDN_flop \out_fifo_reg[7][1][3] (.clk (clk), .d (n_14556), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [3]));
  CDN_flop \out_fifo_reg[7][1][4] (.clk (clk), .d (n_14533), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [4]));
  CDN_flop \out_fifo_reg[7][1][5] (.clk (clk), .d (n_14727), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [5]));
  CDN_flop \out_fifo_reg[7][1][6] (.clk (clk), .d (n_14729), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [6]));
  CDN_flop \out_fifo_reg[7][1][7] (.clk (clk), .d (n_14728), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [7]));
  CDN_flop \out_fifo_reg[7][1][8] (.clk (clk), .d (n_14726), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [8]));
  CDN_flop \out_fifo_reg[7][2][0] (.clk (clk), .d (n_13895), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [0]));
  CDN_flop \out_fifo_reg[7][2][1] (.clk (clk), .d (n_14572), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [1]));
  CDN_flop \out_fifo_reg[7][2][8] (.clk (clk), .d (n_14573), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [8]));
  CDN_flop \out_fifo_reg[7][2][9] (.clk (clk), .d (1'b1), .sena
       (n_13831), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (\out_fifo[7][2] [9]));
  CDN_flop \out_fifo_write_pointer_reg[0] (.clk (clk), .d (n_22039),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[0]));
  CDN_flop \out_fifo_write_pointer_reg[1] (.clk (clk), .d (n_22029),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[1]));
  CDN_flop \out_fifo_write_pointer_reg[2] (.clk (clk), .d (n_22001),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[2]));
  CDN_flop \sh_bit_cnt_reg[0] (.clk (clk), .d (n_13850), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[0]));
  CDN_flop \sh_bit_cnt_reg[1] (.clk (clk), .d (n_22081), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[1]));
  CDN_flop \sh_bit_cnt_reg[2] (.clk (clk), .d (n_22052), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[2]));
  CDN_flop \sh_bit_cnt_reg[3] (.clk (clk), .d (n_14629), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[3]));
  CDN_flop \sh_reg_in_reg[0] (.clk (clk), .d (din), .sena (n_13824),
       .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd (1'b0), .q
       (sh_reg_in[0]));
  CDN_flop \sh_reg_in_reg[1] (.clk (clk), .d (sh_reg_in[0]), .sena
       (n_13824), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (sh_reg_in[1]));
  CDN_flop \sh_reg_in_reg[2] (.clk (clk), .d (sh_reg_in[1]), .sena
       (n_13824), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (sh_reg_in[2]));
  CDN_flop \sh_reg_in_reg[3] (.clk (clk), .d (sh_reg_in[2]), .sena
       (n_13824), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (sh_reg_in[3]));
  CDN_flop \sh_reg_in_reg[4] (.clk (clk), .d (sh_reg_in[3]), .sena
       (n_13824), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (sh_reg_in[4]));
  CDN_flop \sh_reg_in_reg[5] (.clk (clk), .d (sh_reg_in[4]), .sena
       (n_13824), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (sh_reg_in[5]));
  CDN_flop \sh_reg_in_reg[6] (.clk (clk), .d (sh_reg_in[5]), .sena
       (n_13824), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (sh_reg_in[6]));
  CDN_flop \sh_reg_in_reg[7] (.clk (clk), .d (sh_reg_in[6]), .sena
       (n_13824), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (sh_reg_in[7]));
  CDN_flop \sh_reg_in_reg[8] (.clk (clk), .d (sh_reg_in[7]), .sena
       (n_13824), .aclr (1'b0), .apre (1'b0), .srl (n_13823), .srd
       (1'b0), .q (sh_reg_in[8]));
  CDN_flop \sh_reg_out_bit_counter_reg[0] (.clk (clk), .d (n_13909),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[0]));
  CDN_flop \sh_reg_out_bit_counter_reg[1] (.clk (clk), .d (n_22054),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[1]));
  CDN_flop \sh_reg_out_bit_counter_reg[2] (.clk (clk), .d (n_14748),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[2]));
  CDN_flop \sh_reg_out_bit_counter_reg[3] (.clk (clk), .d (n_14750),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[3]));
  CDN_flop \sh_reg_out_bit_counter_reg[4] (.clk (clk), .d (n_14749),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[4]));
  CDN_flop \sh_reg_out_reg[0] (.clk (clk), .d (n_14703), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[0]));
  CDN_flop \sh_reg_out_reg[1] (.clk (clk), .d (n_14764), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[1]));
  CDN_flop \sh_reg_out_reg[2] (.clk (clk), .d (n_14763), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[2]));
  CDN_flop \sh_reg_out_reg[3] (.clk (clk), .d (n_14760), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[3]));
  CDN_flop \sh_reg_out_reg[4] (.clk (clk), .d (n_14759), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[4]));
  CDN_flop \sh_reg_out_reg[5] (.clk (clk), .d (n_14757), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[5]));
  CDN_flop \sh_reg_out_reg[6] (.clk (clk), .d (n_14756), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[6]));
  CDN_flop \sh_reg_out_reg[7] (.clk (clk), .d (n_14754), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[7]));
  CDN_flop \sh_reg_out_reg[8] (.clk (clk), .d (n_14752), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[8]));
  CDN_flop \sh_reg_out_reg[9] (.clk (clk), .d (n_22073), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[9]));
  CDN_flop \sh_reg_out_reg[10] (.clk (clk), .d (n_14765), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[10]));
  CDN_flop \sh_reg_out_reg[11] (.clk (clk), .d (n_14762), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[11]));
  CDN_flop \sh_reg_out_reg[12] (.clk (clk), .d (n_14770), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[12]));
  CDN_flop \sh_reg_out_reg[13] (.clk (clk), .d (n_14766), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[13]));
  CDN_flop \sh_reg_out_reg[14] (.clk (clk), .d (n_14761), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[14]));
  CDN_flop \sh_reg_out_reg[15] (.clk (clk), .d (n_14758), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[15]));
  CDN_flop \sh_reg_out_reg[16] (.clk (clk), .d (n_14753), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[16]));
  CDN_flop \sh_reg_out_reg[17] (.clk (clk), .d (n_14755), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[17]));
  CDN_flop \sh_reg_out_reg[18] (.clk (clk), .d (n_14772), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[18]));
  CDN_flop \sh_reg_out_reg[19] (.clk (clk), .d (n_22061), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[19]));
  CDN_flop \sh_reg_out_reg[20] (.clk (clk), .d (n_14767), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[20]));
  CDN_flop \sh_reg_out_reg[21] (.clk (clk), .d (n_14769), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[21]));
  CDN_flop \sh_reg_out_reg[22] (.clk (clk), .d (n_22060), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[22]));
  CDN_flop \sh_reg_out_reg[23] (.clk (clk), .d (n_22053), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[23]));
  CDN_flop \sh_reg_out_reg[24] (.clk (clk), .d (n_22080), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[24]));
  CDN_flop \sh_reg_out_reg[25] (.clk (clk), .d (n_22079), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[25]));
  CDN_flop \sh_reg_out_reg[26] (.clk (clk), .d (n_22062), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[26]));
  CDN_flop \sh_reg_out_reg[27] (.clk (clk), .d (n_22074), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[27]));
  CDN_flop \sh_reg_out_reg[28] (.clk (clk), .d (n_14768), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[28]));
  CDN_flop \sh_reg_out_reg[29] (.clk (clk), .d (n_14771), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (dout));
endmodule

`ifdef RC_CDN_GENERIC_GATE
`else
module CDN_flop(clk, d, sena, aclr, apre, srl, srd, q);
  input clk, d, sena, aclr, apre, srl, srd;
  output q;
  wire clk, d, sena, aclr, apre, srl, srd;
  wire q;
  reg  qi;
  assign #1 q = qi;
  always 
    @(posedge clk or posedge apre or posedge aclr) 
      if (aclr) 
        qi <= 0;
      else if (apre) 
          qi <= 1;
        else if (srl) 
            qi <= srd;
          else begin
            if (sena) 
              qi <= d;
          end
  initial 
    qi <= 1'b0;
endmodule
`endif
