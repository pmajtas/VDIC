/******************************************************************************
 * (C) Copyright 2022 AGH UST All Rights Reserved
 ******************************************************************************
 * MODULE NAME: vdic_dut_2022
 * VERSION:     1.2
 * DATE:        10-11-2022
 *
 * ABSTRACT:   DUT module for VDIC 2022 labs.
 *              The DUT is RPN calculator type. The arguments are sent first,
 *              than the operator/command.
 *******************************************************************************
 * HISTORY:
 * 20-10-2022 v1.0 Initial version
 * 03-11-2022 v1.1 Added remaining commands
 * 10-11-2022 v1.2 Modifications:
 *            - corrected bug: zero returned for invalid command
 *            - corrected spec: CMD_AND description
 * 
 *******************************************************************************
 * INPUTS
 *    clk      - posedge active clock, always running
 *    rst_n    - synchronous reset active low
 *    din      - serial data input
 *    enable_n - chip enable, active low;

 * OUTPUTS
 *    dout       - serial data output
 *    dout_valid - valid flag for serial data output, active high
 *
 *******************************************************************************

 The clock is always active.
 The DUT operates on the posedge of the clock.
 The DUT receives the data when enable_n is active.
 IMPORTANT: din and dout can operate in parallel - DUT has some internal buffering
 implemented.

 --------------------------------------------------------------------------------
 --- Input data
 --------------------------------------------------------------------------------

 The input data is send serially in WORDs.

 The WORD is always 10 bit long. MSB is sent first.
 The WORD sent to the DUT is either DATA type or CONTROL type.

 DATA = 0bbbbbbbbp
 where:
 - b = 0 or 1, PAYLOAD bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 CONTROL = 1bbbbbbbbp
 where:
 - b = 0 or 1, COMMAND bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 The COMMAND can be:
 00000000 - CMD_NOP, do nothing, remove the data (reset data stack)
 00000001 - CMD_AND, logic AND of the arguments
 00000010 - CMD_OR, logic OR of the arguments
 00000011 - CMD_XOR, logic XOR of the arguments
 00010000 - CMD_ADD, add the arguments
 00100000 - CMD_SUB, subtract other arguments from the first one

 --------------------------------------------------------------------------------
 --- Output data
 --------------------------------------------------------------------------------

 The DUT responds to each CONTROL word, sending 3 WORDS:
 STATUS, DATA, DATA

 STATUS = 1bbbbbbbbp
 where bbbbbbbb is one of:

 00000000 - S_NO_ERROR - data correctly processed
 00000001 - S_MISSING_DATA - missing input data
 00000010 - S_DATA_STACK_OVERFLOW - maximum number of arguments exceeded
 00000100 - S_OUTPUT_FIFO_OVERFLOW - result dropped not possible to process
 00100000 - S_DATA_PARITY_ERROR - input data or command parity error
 01000000 - S_COMMAND_PARITY_ERROR - input data or command parity error
 10000000 - S_INVALID_COMMAND - unknown command detected

 DATA is defined as in the input.
 PAYLOAD of the DATA is 00000000 if the data was NOT processed correctly.

 *******************************************************************************
 * IMPLEMENTATION STATUS
 *******************************************************************************
 *  <Feature>                        <Is implemented>
 *    command CMD_NOP                   YES
 *    command CMD_AND                   YES
 *    command CMD_OR                    YES
 *    command CMD_XOR                   YES
 *    command CMD_ADD                   YES
 *    command CMD_SUB                   YES
 *    status S_NO_ERROR                 YES
 *    status S_MISSING_DATA              NO
 *    status S_DATA_STACK_OVERFLOW       NO
 *    status S_OUTPUT_FIFO_OVERFLOW      NO
 *    status S_DATA_PARITY_ERROR         NO
 *    status S_COMMAND_PARITY_ERROR      NO
 *    status S_INVALID_COMMAND          YES
 *******************************************************************************
 */

module vdic_dut_2022(clk, rst_n, enable_n, din, dout, dout_valid);
  input clk, rst_n, enable_n, din;
  output dout, dout_valid;
  wire clk, rst_n, enable_n, din;
  wire dout, dout_valid;
  wire [7:0] \data_stack_mem[0] ;
  wire [7:0] \data_stack_mem[1] ;
  wire [7:0] \data_stack_mem[2] ;
  wire [7:0] \data_stack_mem[3] ;
  wire [7:0] \data_stack_mem[4] ;
  wire [7:0] \data_stack_mem[5] ;
  wire [7:0] \data_stack_mem[6] ;
  wire [7:0] \data_stack_mem[7] ;
  wire [7:0] \data_stack_mem[8] ;
  wire [3:0] data_stack_pointer;
  wire [2:0] out_fifo_read_pointer;
  wire [2:0] out_fifo_write_pointer;
  wire [3:0] sh_bit_cnt;
  wire [4:0] sh_reg_out_bit_counter;
  wire [9:0] sh_reg_in;
  wire [15:0] result;
  wire [9:0] \out_fifo[4][0] ;
  wire [9:0] \out_fifo[0][0] ;
  wire [9:0] \out_fifo[4][2] ;
  wire [9:0] \out_fifo[0][2] ;
  wire [9:0] \out_fifo[0][1] ;
  wire [9:0] \out_fifo[4][1] ;
  wire [9:0] \out_fifo[6][0] ;
  wire [9:0] \out_fifo[2][2] ;
  wire [9:0] \out_fifo[1][0] ;
  wire [9:0] \out_fifo[5][2] ;
  wire [9:0] \out_fifo[1][2] ;
  wire [9:0] \out_fifo[7][0] ;
  wire [9:0] \out_fifo[5][0] ;
  wire [9:0] \out_fifo[2][0] ;
  wire [9:0] \out_fifo[2][1] ;
  wire [9:0] \out_fifo[3][0] ;
  wire [9:0] \out_fifo[3][1] ;
  wire [9:0] \out_fifo[1][1] ;
  wire [9:0] \out_fifo[7][1] ;
  wire [9:0] \out_fifo[5][1] ;
  wire [9:0] \out_fifo[6][1] ;
  wire [9:0] \out_fifo[6][2] ;
  wire [7:0] status;
  wire [9:0] \out_fifo[3][2] ;
  wire [9:0] \out_fifo[7][2] ;
  wire [29:0] sh_reg_out;
  wire n_11, n_20, n_37, n_100, n_119, n_131, n_139, n_158;
  wire n_168, n_170, n_521, n_523, n_624, n_625, n_633, n_817;
  wire n_827, n_837, n_847, n_857, n_867, n_877, n_887, n_1075;
  wire n_1083, n_1323, n_1325, n_1326, n_1327, n_1329, n_1333, n_1337;
  wire n_1343, n_1345, n_1347, n_1349, n_1351, n_1353, n_1355, n_1357;
  wire n_1359, n_1361, n_1367, n_1371, n_1373, n_1377, n_1379, n_1381;
  wire n_1383, n_1385, n_1387, n_1389, n_1391, n_1393, n_1399, n_1403;
  wire n_1405, n_1409, n_1411, n_1413, n_1415, n_1417, n_1419, n_1421;
  wire n_1423, n_1425, n_1427, n_1429, n_1431, n_1433, n_1435, n_1437;
  wire n_1439, n_1483, n_2033, n_3634, n_3637, n_3649, n_3669, n_3673;
  wire n_3676, n_3683, n_3684, n_3692, n_3693, n_3699, n_3703, n_3710;
  wire n_3711, n_3717, n_3721, n_3726, n_3730, n_3793, n_3902, n_3908;
  wire n_3910, n_4049, n_4050, n_4051, n_4052, n_4053, n_4054, n_4055;
  wire n_4056, n_4081, n_4082, n_4083, n_4084, n_4085, n_4086, n_4087;
  wire n_4088, n_4112, n_4113, n_4114, n_4115, n_4116, n_4117, n_4118;
  wire n_4119, n_4120, n_4144, n_4145, n_4146, n_4147, n_4148, n_4149;
  wire n_4150, n_4151, n_4152, n_4175, n_4176, n_4177, n_4178, n_4179;
  wire n_4180, n_4181, n_4182, n_4183, n_4184, n_4207, n_4208, n_4209;
  wire n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4239;
  wire n_4240, n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248;
  wire n_4330, n_4338, n_4339, n_4340, n_4341, n_4342, n_4343, n_4344;
  wire n_4369, n_4370, n_4371, n_4372, n_4373, n_4374, n_4375, n_4376;
  wire n_4400, n_4401, n_4402, n_4403, n_4404, n_4405, n_4406, n_4407;
  wire n_4408, n_4426, n_4432, n_4433, n_4434, n_4435, n_4436, n_4437;
  wire n_4438, n_4439, n_4440, n_4466, n_4467, n_4468, n_4469, n_4470;
  wire n_4471, n_4472, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500;
  wire n_4501, n_4502, n_4503, n_4504, n_4528, n_4529, n_4530, n_4531;
  wire n_4532, n_4533, n_4534, n_4535, n_4536, n_4615, n_4634, n_4637;
  wire n_4640, n_4642, n_4643, n_4646, n_4684, n_4688, n_4692, n_4696;
  wire n_4700, n_4704, n_4708, n_4712, n_4716, n_4720, n_4724, n_4728;
  wire n_4732, n_4736, n_4740, n_4744, n_4748, n_4752, n_4756, n_4760;
  wire n_4764, n_4768, n_4772, n_4776, n_4780, n_4784, n_4788, n_4792;
  wire n_4796, n_4800, n_4804, n_4808, n_4812, n_4816, n_4820, n_4824;
  wire n_4828, n_4832, n_4836, n_4840, n_4844, n_4848, n_4852, n_4856;
  wire n_4860, n_4864, n_4868, n_4872, n_4876, n_4880, n_4884, n_4888;
  wire n_4892, n_4896, n_4900, n_4904, n_4908, n_4912, n_4916, n_4920;
  wire n_4924, n_4928, n_4932, n_4936, n_4940, n_4944, n_4948, n_4952;
  wire n_4956, n_4960, n_4964, n_4968, n_5004, n_5008, n_5012, n_5016;
  wire n_5019, n_5023, n_5027, n_5031, n_5035, n_5039, n_5043, n_5047;
  wire n_5051, n_5055, n_5059, n_5063, n_5067, n_5071, n_5075, n_5079;
  wire n_5083, n_5087, n_5091, n_5095, n_5099, n_5103, n_5107, n_5111;
  wire n_5115, n_5119, n_5123, n_5127, n_5131, n_5135, n_5139, n_5143;
  wire n_5147, n_5151, n_5155, n_5159, n_5163, n_5167, n_5171, n_5175;
  wire n_5179, n_5183, n_5187, n_5191, n_5195, n_5199, n_5203, n_5207;
  wire n_5211, n_5215, n_5219, n_5223, n_5227, n_5231, n_5235, n_5239;
  wire n_5243, n_5247, n_5251, n_5255, n_5259, n_5263, n_5267, n_5271;
  wire n_5275, n_5279, n_5283, n_5287, n_5291, n_5295, n_5299, n_5303;
  wire n_5307, n_5311, n_5315, n_5319, n_5323, n_5327, n_5331, n_5335;
  wire n_5339, n_5343, n_5347, n_5351, n_5355, n_5359, n_5363, n_5367;
  wire n_5371, n_5375, n_5379, n_5383, n_5387, n_5391, n_5395, n_5399;
  wire n_5403, n_5407, n_5411, n_5415, n_5419, n_5423, n_5427, n_5431;
  wire n_5435, n_5439, n_5443, n_5447, n_5451, n_5455, n_5459, n_5463;
  wire n_5467, n_5471, n_5475, n_5479, n_5483, n_5487, n_5491, n_5495;
  wire n_5499, n_5503, n_5507, n_5511, n_5515, n_5519, n_5523, n_5527;
  wire n_5531, n_5535, n_5539, n_5543, n_5547, n_5551, n_5555, n_5559;
  wire n_5563, n_5567, n_5571, n_5575, n_5579, n_5583, n_5587, n_5591;
  wire n_5595, n_5599, n_5603, n_5607, n_5611, n_5615, n_5619, n_5622;
  wire n_5625, n_5628, n_5631, n_5635, n_5643, n_5647, n_5651, n_5653;
  wire n_5655, n_5657, n_5659, n_5661, n_5663, n_5665, n_5667, n_5669;
  wire n_5673, n_5675, n_5677, n_5679, n_5681, n_5683, n_5685, n_5687;
  wire n_5689, n_5693, n_5695, n_5709, n_5711, n_5715, n_5719, n_5723;
  wire n_5727, n_5731, n_5735, n_5739, n_5743, n_5747, n_5751, n_5755;
  wire n_5759, n_5763, n_5767, n_5771, n_5775, n_5779, n_5783, n_5787;
  wire n_5791, n_5795, n_5799, n_5803, n_5807, n_11305, n_11312,
       n_11318;
  wire n_11331, n_11358, n_11432, n_11449, n_11474, n_11478, n_11480,
       n_11483;
  wire n_11521, n_11540, n_11572, n_11576, n_11578, n_11581, n_11622,
       n_11641;
  wire n_11673, n_11677, n_11679, n_11682, n_11723, n_11742, n_11774,
       n_11778;
  wire n_11780, n_11783, n_11824, n_11843, n_11875, n_11879, n_11881,
       n_11884;
  wire n_11925, n_11944, n_11973, n_11974, n_11976, n_11978, n_11980,
       n_11982;
  wire n_11985, n_11986, n_12027, n_12045, n_12070, n_12074, n_12076,
       n_12079;
  wire n_12119, n_12141, n_12166, n_12170, n_12172, n_12175, n_12218,
       n_12240;
  wire n_12265, n_12269, n_12271, n_12274, n_12317, n_12339, n_12364,
       n_12368;
  wire n_12370, n_12373, n_12416, n_12438, n_12463, n_12467, n_12469,
       n_12472;
  wire n_12515, n_12537, n_12553, n_12562, n_12563, n_12566, n_12567,
       n_12568;
  wire n_12569, n_12571, n_12606, n_12622, n_12639, n_12643, n_12645,
       n_12648;
  wire n_12683, n_12699, n_12716, n_12720, n_12722, n_12725, n_12732,
       n_12733;
  wire n_12734, n_12738, n_12739, n_12753, n_12754, n_12755, n_12756,
       n_12757;
  wire n_12758, n_12759, n_12760, n_12761, n_12762, n_12764, n_12765,
       n_12766;
  wire n_12767, n_12768, n_12769, n_12772, n_12774, n_12775, n_12777,
       n_12779;
  wire n_12780, n_12782, n_12785, n_12786, n_12801, n_12803, n_12806,
       n_12808;
  wire n_12809, n_12813, n_12814, n_12824, n_12827, n_12847, n_12853,
       n_12854;
  wire n_12860, n_12861, n_12862, n_12863, n_12864, n_12866, n_12869,
       n_12870;
  wire n_12871, n_12872, n_12895, n_12896, n_12897, n_12898, n_12904,
       n_12905;
  wire n_12917, n_12920, n_12921, n_12929, n_12932, n_12933, n_12941,
       n_13105;
  wire n_13106, n_13107, n_13108, n_13109, n_13110, n_13111, n_13121,
       n_13123;
  wire n_13131, n_13134, n_13135, n_13137, n_13138, n_13139, n_13140,
       n_13141;
  wire n_13142, n_13146, n_13147, n_13183, n_13189, n_13190, n_13191,
       n_13197;
  wire n_13203, n_13214, n_13215, n_13220, n_13233, n_13242, n_13244,
       n_13400;
  wire n_13401, n_13402, n_13403, n_13404, n_13405, n_13406, n_13407,
       n_13409;
  wire n_13428, n_13439, n_13443, n_13449, n_13450, n_13452, n_13533,
       n_13536;
  wire n_13538, n_13608, n_13744, n_13764, n_13765, n_13766, n_13767,
       n_13768;
  wire n_13769, n_13770, n_13772, n_13773, n_13774, n_13775, n_13776,
       n_13777;
  wire n_13778, n_13779, n_13780, n_13781, n_13782, n_13783, n_13784,
       n_13785;
  wire n_13788, n_13789, n_13791, n_13792, n_13793, n_13794, n_13795,
       n_13797;
  wire n_13798, n_13803, n_13804, n_13805, n_13806, n_13807, n_13808,
       n_13809;
  wire n_13811, n_13812, n_13813, n_13814, n_13815, n_13816, n_13817,
       n_13818;
  wire n_13821, n_13822, n_13825, n_13826, n_13827, n_13828, n_13830,
       n_13831;
  wire n_13832, n_13898, n_13900, n_13901, n_13902, n_13903, n_13904,
       n_13905;
  wire n_13906, n_13907, n_13908, n_13909, n_13911, n_13912, n_13913,
       n_13914;
  wire n_13915, n_13916, n_13917, n_13918, n_13919, n_13920, n_13921,
       n_13922;
  wire n_13925, n_13928, n_13931, n_13932, n_13933, n_13934, n_13935,
       n_13936;
  wire n_13938, n_13939, n_13940, n_13941, n_13942, n_13943, n_13944,
       n_13945;
  wire n_13946, n_13947, n_13948, n_13949, n_13950, n_13951, n_13952,
       n_13953;
  wire n_13956, n_13957, n_13958, n_13959, n_13960, n_13961, n_13962,
       n_13964;
  wire n_13965, n_13966, n_13967, n_13969, n_13970, n_13971, n_13972,
       n_13975;
  wire n_13976, n_13977, n_13978, n_13979, n_13980, n_13981, n_13982,
       n_13983;
  wire n_13984, n_13985, n_13986, n_13987, n_13988, n_13989, n_13990,
       n_13991;
  wire n_13992, n_13993, n_13994, n_13995, n_13996, n_13998, n_14000,
       n_14003;
  wire n_14009, n_14010, n_14011, n_14012, n_14013, n_14014, n_14016,
       n_14023;
  wire n_14024, n_14025, n_14029, n_14030, n_14031, n_14032, n_14034,
       n_14035;
  wire n_14036, n_14038, n_14039, n_14040, n_14041, n_14043, n_14045,
       n_14047;
  wire n_14049, n_14051, n_14052, n_14053, n_14054, n_14055, n_14056,
       n_14058;
  wire n_14060, n_14063, n_14064, n_14069, n_14070, n_14072, n_14075,
       n_14076;
  wire n_14078, n_14084, n_14085, n_14086, n_14087, n_14089, n_14090,
       n_14093;
  wire n_14096, n_14098, n_14099, n_14100, n_14102, n_14103, n_14107,
       n_14108;
  wire n_14109, n_14110, n_14111, n_14112, n_14113, n_14114, n_14116,
       n_14120;
  wire n_14125, n_14126, n_14127, n_14128, n_14130, n_14131, n_14132,
       n_14133;
  wire n_14134, n_14135, n_14136, n_14137, n_14140, n_14141, n_14142,
       n_14143;
  wire n_14144, n_14145, n_14147, n_14148, n_14150, n_14151, n_14152,
       n_14153;
  wire n_14159, n_14160, n_14163, n_14164, n_14165, n_14166, n_14167,
       n_14168;
  wire n_14170, n_14171, n_14172, n_14173, n_14174, n_14175, n_14178,
       n_14180;
  wire n_14181, n_14184, n_14189, n_14190, n_14191, n_14192, n_14193,
       n_14194;
  wire n_14195, n_14196, n_14197, n_14198, n_14199, n_14200, n_14201,
       n_14202;
  wire n_14203, n_14204, n_14205, n_14206, n_14207, n_14208, n_14209,
       n_14210;
  wire n_14211, n_14212, n_14213, n_14214, n_14215, n_14216, n_14217,
       n_14218;
  wire n_14219, n_14220, n_14221, n_14222, n_14223, n_14224, n_14225,
       n_14226;
  wire n_14227, n_14228, n_14229, n_14230, n_14231, n_14232, n_14233,
       n_14234;
  wire n_14236, n_14237, n_14238, n_14240, n_14242, n_14243, n_14244,
       n_14246;
  wire n_14247, n_14248, n_14249, n_14250, n_14252, n_14253, n_14254,
       n_14255;
  wire n_14256, n_14257, n_14258, n_14259, n_14260, n_14261, n_14262,
       n_14263;
  wire n_14264, n_14265, n_14266, n_14267, n_14268, n_14269, n_14270,
       n_14271;
  wire n_14272, n_14273, n_14274, n_14275, n_14276, n_14277, n_14278,
       n_14279;
  wire n_14280, n_14281, n_14282, n_14283, n_14284, n_14286, n_14287,
       n_14288;
  wire n_14289, n_14290, n_14291, n_14292, n_14293, n_14294, n_14295,
       n_14296;
  wire n_14297, n_14298, n_14299, n_14300, n_14301, n_14302, n_14303,
       n_14304;
  wire n_14305, n_14307, n_14308, n_14309, n_14310, n_14311, n_14312,
       n_14313;
  wire n_14314, n_14315, n_14316, n_14317, n_14463, n_14464, n_14465,
       n_14466;
  wire n_14467, n_14468, n_14469, n_14470, n_14471, n_14472, n_14473,
       n_14475;
  wire n_14477, n_14479, n_14480, n_14482, n_14483, n_14485, n_14487,
       n_14489;
  wire n_14491, n_14493, n_14494, n_14495, n_14496, n_14497, n_14499,
       n_14500;
  wire n_14501, n_14502, n_14504, n_14505, n_14506, n_14509, n_14510,
       n_14512;
  wire n_14513, n_14514, n_14515, n_14516, n_14517, n_14518, n_14519,
       n_14520;
  wire n_14521, n_14523, n_14524, n_14526, n_14527, n_14529, n_14530,
       n_14532;
  wire n_14533, n_14534, n_14535, n_14536, n_14537, n_14538, n_14539,
       n_14540;
  wire n_14544, n_14545, n_14546, n_14549, n_14550, n_14551, n_14552,
       n_14553;
  wire n_14554, n_14556, n_14557, n_14558, n_14559, n_14566, n_14567,
       n_14569;
  wire n_14570, n_14571, n_14572, n_14574, n_14575, n_14576, n_14578,
       n_14580;
  wire n_14581, n_14582, n_14583, n_14584, n_14585, n_14586, n_14587,
       n_14588;
  wire n_14589, n_14590, n_14591, n_14592, n_14593, n_14594, n_14621,
       n_14622;
  wire n_14623, n_14624, n_14625, n_14626, n_14627, n_14628, n_14635,
       n_14636;
  wire n_14637, n_14642, n_14643, n_14648, n_14649, n_14654, n_14655,
       n_14658;
  wire n_14661, n_14664, n_14667, n_14670, n_14673, n_14676, n_14681,
       n_14682;
  wire n_14685, n_14688, n_14697, n_14698, n_14699, n_14700, n_14705,
       n_14706;
  wire n_14717, n_14718, n_14721, n_14730, n_14731, n_14732, n_14733,
       n_14740;
  wire n_14741, n_14742, n_14745, n_14748, n_14751, n_14754, n_14757,
       n_14764;
  wire n_14765, n_14766, n_14795, n_14796, n_14797, n_14798, n_14799,
       n_14800;
  wire n_14801, n_14802, n_14803, n_14804, n_14805, n_14806, n_14807,
       n_14808;
  wire n_14811, n_14814, n_14817, n_14820, n_14823, n_14826, n_14833,
       n_14834;
  wire n_14835, n_14862, n_14863, n_14864, n_14865, n_14866, n_14867,
       n_14868;
  wire n_14869, n_14870, n_14871, n_14872, n_14873, n_14874, n_14901,
       n_14902;
  wire n_14903, n_14904, n_14905, n_14906, n_14907, n_14908, n_14909,
       n_14910;
  wire n_14911, n_14912, n_14913, n_14916, n_14919, n_14922, n_14925,
       n_14934;
  wire n_14935, n_14936, n_14937, n_14946, n_14947, n_14948, n_14949,
       n_14958;
  wire n_14959, n_14960, n_14961, n_14968, n_14969, n_14970, n_14975,
       n_14976;
  wire n_14985, n_14986, n_14987, n_14988, n_14995, n_14996, n_14997,
       n_15000;
  wire n_15015, n_15016, n_15017, n_15018, n_15019, n_15020, n_15021,
       n_15034;
  wire n_15035, n_15036, n_15037, n_15038, n_15039, n_15064, n_15065,
       n_15066;
  wire n_15067, n_15068, n_15069, n_15070, n_15071, n_15072, n_15073,
       n_15074;
  wire n_15075, n_15088, n_15089, n_15090, n_15091, n_15092, n_15093,
       n_15106;
  wire n_15107, n_15108, n_15109, n_15110, n_15111, n_15130, n_15131,
       n_15132;
  wire n_15133, n_15134, n_15135, n_15144, n_15145, n_15146, n_15147,
       n_15156;
  wire n_15157, n_15158, n_15159, n_15186, n_15187, n_15188, n_15189,
       n_15190;
  wire n_15191, n_15192, n_15193, n_15194, n_15195, n_15196, n_15197,
       n_15198;
  wire n_15207, n_15208, n_15209, n_15210, n_15239, n_15240, n_15241,
       n_15242;
  wire n_15243, n_15244, n_15245, n_15246, n_15247, n_15248, n_15249,
       n_15250;
  wire n_15251, n_15252, n_15261, n_15262, n_15263, n_15264, n_15273,
       n_15274;
  wire n_15275, n_15276, n_15279, n_15282, n_15285, n_15288, n_15299,
       n_15300;
  wire n_15305, n_15306, n_15309, n_15316, n_15317, n_15318, n_15321,
       n_15326;
  wire n_15327, n_15330, n_15333, n_15336, n_15339, n_15342, n_15363,
       n_15364;
  wire n_15365, n_15366, n_15367, n_15368, n_15369, n_15370, n_15371,
       n_15372;
  wire n_15375, n_15384, n_15385, n_15386, n_15387, n_15390, n_15393,
       n_15418;
  wire n_15419, n_15420, n_15421, n_15422, n_15423, n_15424, n_15425,
       n_15426;
  wire n_15427, n_15428, n_15429, n_15434, n_15435, n_15440, n_15441,
       n_15446;
  wire n_15447, n_15452, n_15453, n_15456, n_15463, n_15464, n_15465,
       n_15472;
  wire n_15473, n_15474, n_15479, n_15480, n_15483, n_15486, n_15489,
       n_15494;
  wire n_15495, n_15498, n_15501, n_15504, n_15507, n_15514, n_15515,
       n_15516;
  wire n_15521, n_15522, n_15527, n_15536, n_15537, n_15542, n_15543,
       n_15554;
  wire n_15555, n_15556, n_15558, n_15564, n_15567, n_15576, n_15577,
       n_15578;
  wire n_15579, n_15588, n_15589, n_15590, n_15591, n_15594, n_15597,
       n_15600;
  wire n_15605, n_15606, n_15617, n_15618, n_15619, n_15620, n_15621,
       n_15624;
  wire n_15629, n_15630, n_15633, n_15638, n_15639, n_15644, n_15645,
       n_15648;
  wire n_15653, n_15654, n_15659, n_15660, n_15665, n_15666, n_15671,
       n_15672;
  wire n_15677, n_15678, n_15683, n_15684, n_15689, n_15690, n_15695,
       n_15696;
  wire n_15701, n_15702, n_15707, n_15708, n_15713, n_15714, n_15719,
       n_15720;
  wire n_15725, n_15726, n_15731, n_15732, n_15737, n_15738, n_15743,
       n_15744;
  wire n_15749, n_15750, n_15755, n_15756, n_15761, n_15762, n_15767,
       n_15768;
  wire n_15773, n_15774, n_15779, n_15780, n_15785, n_15786, n_15791,
       n_15792;
  wire n_15797, n_15798, n_15803, n_15804, n_15809, n_15810, n_15815,
       n_15816;
  wire n_15821, n_15822, n_15827, n_15828, n_15833, n_15834, n_15839,
       n_15840;
  wire n_15845, n_15846, n_15851, n_15852, n_15857, n_15858, n_15863,
       n_15864;
  wire n_15869, n_15870, n_15875, n_15876, n_15881, n_15882, n_15887,
       n_15888;
  wire n_15893, n_15894, n_15899, n_15900, n_15905, n_15906, n_15911,
       n_15912;
  wire n_15917, n_15918, n_15923, n_15924, n_15929, n_15930, n_15935,
       n_15936;
  wire n_15943, n_15944, n_15945, n_15950, n_15951, n_15954, n_15957,
       n_15960;
  wire n_15965, n_15966, n_15973, n_15974, n_15975, n_15982, n_15983,
       n_15984;
  wire n_15989, n_15990, n_15993, n_15996, n_16001, n_16002, n_16007,
       n_16008;
  wire n_16013, n_16014, n_16019, n_16020, n_16025, n_16026, n_16031,
       n_16032;
  wire n_16037, n_16038, n_16043, n_16044, n_16049, n_16050, n_16055,
       n_16056;
  wire n_16061, n_16062, n_16067, n_16068, n_16073, n_16074, n_16079,
       n_16080;
  wire n_16085, n_16086, n_16091, n_16092, n_16097, n_16098, n_16103,
       n_16104;
  wire n_16109, n_16110, n_16115, n_16116, n_16121, n_16122, n_16127,
       n_16128;
  wire n_16133, n_16134, n_16139, n_16140, n_16145, n_16146, n_16151,
       n_16152;
  wire n_16157, n_16158, n_16163, n_16164, n_16169, n_16170, n_16175,
       n_16176;
  wire n_16181, n_16182, n_16187, n_16188, n_16193, n_16194, n_16199,
       n_16200;
  wire n_16205, n_16206, n_16211, n_16212, n_16217, n_16218, n_16223,
       n_16224;
  wire n_16253, n_16254, n_16255, n_16256, n_16257, n_16258, n_16259,
       n_16260;
  wire n_16261, n_16262, n_16263, n_16264, n_16265, n_16266, n_16271,
       n_16272;
  wire n_16277, n_16278, n_16283, n_16284, n_16289, n_16290, n_16323,
       n_16324;
  wire n_16325, n_16326, n_16327, n_16328, n_16329, n_16330, n_16331,
       n_16332;
  wire n_16333, n_16334, n_16335, n_16336, n_16337, n_16338, n_16371,
       n_16372;
  wire n_16373, n_16374, n_16375, n_16376, n_16377, n_16378, n_16379,
       n_16380;
  wire n_16381, n_16382, n_16383, n_16384, n_16385, n_16386, n_16419,
       n_16420;
  wire n_16421, n_16422, n_16423, n_16424, n_16425, n_16426, n_16427,
       n_16428;
  wire n_16429, n_16430, n_16431, n_16432, n_16433, n_16434, n_16467,
       n_16468;
  wire n_16469, n_16470, n_16471, n_16472, n_16473, n_16474, n_16475,
       n_16476;
  wire n_16477, n_16478, n_16479, n_16480, n_16481, n_16482, n_16515,
       n_16516;
  wire n_16517, n_16518, n_16519, n_16520, n_16521, n_16522, n_16523,
       n_16524;
  wire n_16525, n_16526, n_16527, n_16528, n_16529, n_16530, n_16563,
       n_16564;
  wire n_16565, n_16566, n_16567, n_16568, n_16569, n_16570, n_16571,
       n_16572;
  wire n_16573, n_16574, n_16575, n_16576, n_16577, n_16578, n_16611,
       n_16612;
  wire n_16613, n_16614, n_16615, n_16616, n_16617, n_16618, n_16619,
       n_16620;
  wire n_16621, n_16622, n_16623, n_16624, n_16625, n_16626, n_16659,
       n_16660;
  wire n_16661, n_16662, n_16663, n_16664, n_16665, n_16666, n_16667,
       n_16668;
  wire n_16669, n_16670, n_16671, n_16672, n_16673, n_16674, n_16707,
       n_16708;
  wire n_16709, n_16710, n_16711, n_16712, n_16713, n_16714, n_16715,
       n_16716;
  wire n_16717, n_16718, n_16719, n_16720, n_16721, n_16722, n_16755,
       n_16756;
  wire n_16757, n_16758, n_16759, n_16760, n_16761, n_16762, n_16763,
       n_16764;
  wire n_16765, n_16766, n_16767, n_16768, n_16769, n_16770, n_16803,
       n_16804;
  wire n_16805, n_16806, n_16807, n_16808, n_16809, n_16810, n_16811,
       n_16812;
  wire n_16813, n_16814, n_16815, n_16816, n_16817, n_16818, n_16851,
       n_16852;
  wire n_16853, n_16854, n_16855, n_16856, n_16857, n_16858, n_16859,
       n_16860;
  wire n_16861, n_16862, n_16863, n_16864, n_16865, n_16866, n_16899,
       n_16900;
  wire n_16901, n_16902, n_16903, n_16904, n_16905, n_16906, n_16907,
       n_16908;
  wire n_16909, n_16910, n_16911, n_16912, n_16913, n_16914, n_16947,
       n_16948;
  wire n_16949, n_16950, n_16951, n_16952, n_16953, n_16954, n_16955,
       n_16956;
  wire n_16957, n_16958, n_16959, n_16960, n_16961, n_16962, n_16995,
       n_16996;
  wire n_16997, n_16998, n_16999, n_17000, n_17001, n_17002, n_17003,
       n_17004;
  wire n_17005, n_17006, n_17007, n_17008, n_17009, n_17010, n_17043,
       n_17044;
  wire n_17045, n_17046, n_17047, n_17048, n_17049, n_17050, n_17051,
       n_17052;
  wire n_17053, n_17054, n_17055, n_17056, n_17057, n_17058, n_17091,
       n_17092;
  wire n_17093, n_17094, n_17095, n_17096, n_17097, n_17098, n_17099,
       n_17100;
  wire n_17101, n_17102, n_17103, n_17104, n_17105, n_17106, n_17139,
       n_17140;
  wire n_17141, n_17142, n_17143, n_17144, n_17145, n_17146, n_17147,
       n_17148;
  wire n_17149, n_17150, n_17151, n_17152, n_17153, n_17154, n_17187,
       n_17188;
  wire n_17189, n_17190, n_17191, n_17192, n_17193, n_17194, n_17195,
       n_17196;
  wire n_17197, n_17198, n_17199, n_17200, n_17201, n_17202, n_17235,
       n_17236;
  wire n_17237, n_17238, n_17239, n_17240, n_17241, n_17242, n_17243,
       n_17244;
  wire n_17245, n_17246, n_17247, n_17248, n_17249, n_17250, n_17283,
       n_17284;
  wire n_17285, n_17286, n_17287, n_17288, n_17289, n_17290, n_17291,
       n_17292;
  wire n_17293, n_17294, n_17295, n_17296, n_17297, n_17298, n_17303,
       n_17304;
  wire n_17309, n_17310, n_17315, n_17319, n_17324, n_17325, n_17330,
       n_17331;
  wire n_17336, n_17337, n_17342, n_17343, n_17348, n_17349, n_17354,
       n_17355;
  wire n_17366, n_17367, n_17368, n_17369, n_17370, n_17375, n_17376,
       n_17383;
  wire n_17384, n_17385, n_17390, n_17391, n_17398, n_17399, n_17400,
       n_17405;
  wire n_17406, n_17411, n_17412, n_17417, n_17418, n_17423, n_17424,
       n_17429;
  wire n_17430, n_17435, n_17441, n_17453, n_17454, n_17455, n_17456,
       n_17457;
  wire n_17462, n_17463, n_17474, n_17475, n_17476, n_17477, n_17478,
       n_17483;
  wire n_17484, n_17489, n_17490, n_17495, n_17496, n_17501, n_17502,
       n_17507;
  wire n_17508, n_17513, n_17514, n_17519, n_17520, n_17525, n_17526,
       n_17531;
  wire n_17532, n_17537, n_17538, n_17543, n_17544, n_17549, n_17550,
       n_17555;
  wire n_17556, n_17561, n_17562, n_17567, n_17568, n_17573, n_17574,
       n_17579;
  wire n_17580, n_17585, n_17586, n_17591, n_17592, n_17597, n_17598,
       n_17603;
  wire n_17604, n_17609, n_17610, n_17615, n_17621, n_17622, n_17627,
       n_17633;
  wire n_17639, n_17647, n_17648, n_17649, n_17654, n_17655, n_17660,
       n_17661;
  wire n_17666, n_17667, n_17672, n_17673, n_17678, n_17679, n_17684,
       n_17685;
  wire n_17690, n_17691, n_17696, n_17697, n_17702, n_17703, n_17708,
       n_17709;
  wire n_17714, n_17715, n_17720, n_17721, n_17726, n_17727, n_17732,
       n_17738;
  wire n_17739, n_17744, n_17745, n_17750, n_17751, n_17756, n_17757,
       n_17762;
  wire n_17763, n_17766, n_17769, n_17774, n_17775, n_17780, n_17781,
       n_17792;
  wire n_17793, n_17794, n_17795, n_17796, n_17801, n_17802, n_17807,
       n_17808;
  wire n_17813, n_17814, n_17819, n_17820, n_17825, n_17826, n_17831,
       n_17832;
  wire n_17837, n_17838, n_17843, n_17847, n_17856, n_17857, n_17858,
       n_17859;
  wire n_17862, n_17865, n_17870, n_17871, n_17876, n_17877, n_17882,
       n_17883;
  wire n_17886, n_17891, n_17897, n_17898, n_17905, n_17906, n_17907,
       n_17910;
  wire n_17915, n_17916, n_17921, n_17922, n_17927, n_17928, n_17933,
       n_17934;
  wire n_17939, n_17940, n_17945, n_17946, n_17951, n_17952, n_17957,
       n_17958;
  wire n_17963, n_17964, n_17969, n_17970, n_17975, n_17976, n_17981,
       n_17982;
  wire n_17987, n_17988, n_17993, n_17994, n_17999, n_18000, n_18003,
       n_18006;
  wire n_18011, n_18012, n_18017, n_18018, n_18023, n_18024, n_18029,
       n_18030;
  wire n_18035, n_18036, n_18043, n_18044, n_18045, n_18048, n_18053,
       n_18054;
  wire n_18057, n_18060, n_18065, n_18066, n_18071, n_18072, n_18077,
       n_18078;
  wire n_18083, n_18084, n_18089, n_18090, n_18093, n_18096, n_18101,
       n_18102;
  wire n_18121, n_18122, n_18123, n_18124, n_18125, n_18126, n_18127,
       n_18128;
  wire n_18129, n_18134, n_18135, n_18140, n_18141, n_18146, n_18147,
       n_18152;
  wire n_18153, n_18158, n_18159, n_18164, n_18165, n_18170, n_18171,
       n_18176;
  wire n_18177, n_18182, n_18183, n_18186, n_18191, n_18195, n_18198,
       n_18201;
  wire n_18206, n_18207, n_18218, n_18219, n_18220, n_18221, n_18222,
       n_18227;
  wire n_18228, n_18233, n_18234, n_18237, n_18240, n_18243, n_18248,
       n_18249;
  wire n_18256, n_18257, n_18258, n_18263, n_18264, n_18269, n_18270,
       n_18275;
  wire n_18276, n_18279, n_18282, n_18287, n_18288, n_18291, n_18294,
       n_18313;
  wire n_18314, n_18315, n_18316, n_18317, n_18318, n_18319, n_18320,
       n_18321;
  wire n_18326, n_18327, n_18332, n_18333, n_18338, n_18339, n_18344,
       n_18345;
  wire n_18350, n_18351, n_18356, n_18357, n_18362, n_18363, n_18368,
       n_18369;
  wire n_18372, n_18379, n_18380, n_18381, n_18384, n_18387, n_18392,
       n_18393;
  wire n_18398, n_18399, n_18402, n_18405, n_18424, n_18425, n_18426,
       n_18427;
  wire n_18428, n_18429, n_18430, n_18431, n_18432, n_18437, n_18438,
       n_18443;
  wire n_18444, n_18449, n_18450, n_18455, n_18456, n_18461, n_18462,
       n_18467;
  wire n_18468, n_18473, n_18474, n_18479, n_18480, n_18485, n_18486,
       n_18489;
  wire n_18494, n_18495, n_18500, n_18501, n_18504, n_18507, n_18510,
       n_18517;
  wire n_18518, n_18519, n_18522, n_18527, n_18528, n_18531, n_18550,
       n_18551;
  wire n_18552, n_18553, n_18554, n_18555, n_18556, n_18557, n_18558,
       n_18563;
  wire n_18564, n_18569, n_18570, n_18575, n_18576, n_18581, n_18582,
       n_18587;
  wire n_18588, n_18593, n_18594, n_18599, n_18600, n_18605, n_18606,
       n_18611;
  wire n_18612, n_18615, n_18620, n_18621, n_18626, n_18627, n_18632,
       n_18633;
  wire n_18640, n_18641, n_18642, n_18645, n_18648, n_18667, n_18668,
       n_18669;
  wire n_18670, n_18671, n_18672, n_18673, n_18674, n_18675, n_18680,
       n_18681;
  wire n_18686, n_18687, n_18692, n_18693, n_18698, n_18699, n_18704,
       n_18705;
  wire n_18710, n_18711, n_18716, n_18717, n_18722, n_18723, n_18726,
       n_18729;
  wire n_18732, n_18737, n_18738, n_18745, n_18746, n_18747, n_18750,
       n_18758;
  wire n_18759, n_18778, n_18779, n_18780, n_18781, n_18782, n_18783,
       n_18784;
  wire n_18785, n_18786, n_18791, n_18792, n_18797, n_18798, n_18803,
       n_18804;
  wire n_18809, n_18810, n_18815, n_18816, n_18821, n_18822, n_18827,
       n_18828;
  wire n_18833, n_18834, n_18839, n_18840, n_18843, n_18846, n_18849,
       n_18852;
  wire n_18857, n_18858, n_18861, n_18866, n_18867, n_18872, n_18873,
       n_18878;
  wire n_18879, n_18884, n_18885, n_18890, n_18891, n_18896, n_18897,
       n_18902;
  wire n_18903, n_18906, n_18909, n_18912, n_18915, n_18918, n_18921,
       n_18924;
  wire n_18927, n_18930, n_18933, n_18936, n_18939, n_18942, n_18945,
       n_18948;
  wire n_18951, n_18954, n_18957, n_18960, n_18963, n_18966, n_18969,
       n_18972;
  wire n_18975, n_18978, n_18981, n_18984, n_18987, n_18990, n_18993,
       n_18996;
  wire n_18999, n_19004, n_19005, n_19010, n_19011, n_19018, n_19019,
       n_19020;
  wire n_19039, n_19040, n_19041, n_19042, n_19043, n_19044, n_19045,
       n_19046;
  wire n_19047, n_19052, n_19053, n_19058, n_19059, n_19064, n_19065,
       n_19070;
  wire n_19071, n_19076, n_19077, n_19082, n_19083, n_19088, n_19089,
       n_19094;
  wire n_19095, n_19100, n_19101, n_19106, n_19107, n_19112, n_19113,
       n_19118;
  wire n_19119, n_19124, n_19125, n_19130, n_19131, n_19136, n_19137,
       n_19142;
  wire n_19143, n_19148, n_19149, n_19154, n_19155, n_19160, n_19161,
       n_19166;
  wire n_19167, n_19172, n_19173, n_19178, n_19179, n_19184, n_19185,
       n_19190;
  wire n_19191, n_19196, n_19197, n_19202, n_19203, n_19208, n_19209,
       n_19214;
  wire n_19215, n_19220, n_19221, n_19226, n_19227, n_19232, n_19233,
       n_19238;
  wire n_19239, n_19244, n_19245, n_19250, n_19251, n_19256, n_19257,
       n_19262;
  wire n_19263, n_19268, n_19269, n_19274, n_19275, n_19280, n_19281,
       n_19286;
  wire n_19287, n_19292, n_19293, n_19298, n_19299, n_19304, n_19305,
       n_19310;
  wire n_19311, n_19316, n_19317, n_19322, n_19323, n_19328, n_19329,
       n_19334;
  wire n_19335, n_19340, n_19341, n_19344, n_19347, n_19350, n_19353,
       n_19356;
  wire n_19361, n_19362, n_19365, n_19368, n_19371, n_19374, n_19377,
       n_19380;
  wire n_19383, n_19386, n_19389, n_19392, n_19395, n_19398, n_19401,
       n_19404;
  wire n_19407, n_19410, n_19413, n_19416, n_19419, n_19422, n_19425,
       n_19428;
  wire n_19431, n_19434, n_19437, n_19440, n_19443, n_19446, n_19449,
       n_19452;
  wire n_19455, n_19458, n_19461, n_19464, n_19467, n_19470, n_19473,
       n_19476;
  wire n_19479, n_19482, n_19485, n_19488, n_19491, n_19494, n_19497,
       n_19500;
  wire n_19503, n_19506, n_19509, n_19512, n_19515, n_19518, n_19521,
       n_19524;
  wire n_19527, n_19530, n_19533, n_19536, n_19539, n_19542, n_19545,
       n_19548;
  wire n_19551, n_19554, n_19557, n_19560, n_19563, n_19566, n_19569,
       n_19572;
  wire n_19575, n_19578, n_19581, n_19584, n_19587, n_19590, n_19593,
       n_19596;
  wire n_19601, n_19602, n_19609, n_19610, n_19611, n_20604, n_20605,
       n_20606;
  wire n_20607, n_20608, n_20609, n_20612, n_20613, n_20614, n_20615,
       n_20616;
  wire n_20617, n_20618, n_20619, n_20620, n_20621, n_20622, n_20623,
       n_20624;
  wire n_20625, n_20626, n_20627, n_20628, n_20629, n_20632, n_20633,
       n_20634;
  wire n_20635, n_20636, n_20637, n_20638, n_20639, n_20642, n_20643,
       n_20644;
  wire n_20645, n_20646, n_20647, n_20648, n_20649, n_20652, n_20653,
       n_20654;
  wire n_20655, n_20656, n_20657, n_20658, n_20659, n_20660, n_20661,
       n_20662;
  wire n_20663, n_20664, n_20665, n_20668, n_20669, n_20670, n_20671,
       n_20672;
  wire n_20673, n_20674, n_20675, n_20676, n_20677, n_20678, n_20679,
       n_20680;
  wire n_20681, n_20682, n_20683, n_20684, n_20685, n_20686, n_20687,
       n_20688;
  wire n_20689, n_20690, n_20691, n_20692, n_20693, n_20694, n_20695,
       n_20696;
  wire n_20697, n_20698, n_20699, n_20700, n_20701, n_20702, n_20703,
       n_20704;
  wire n_20705, n_20706, n_20707, n_20710, n_20711, n_20712, n_20713,
       n_20714;
  wire n_20715, n_20716, n_20717, n_20718, n_20719, n_20720, n_20721,
       n_20722;
  wire n_20723, n_20724, n_20725, n_20726, n_20727, n_20728, n_20729,
       n_20730;
  wire n_20731, n_20732, n_20733, n_20734, n_20735, n_20736, n_20737,
       n_20738;
  wire n_20739, n_20740, n_20741, n_20742, n_20743, n_20744, n_20745,
       n_20746;
  wire n_20747, n_20748, n_20749, n_20750, n_20751, n_20752, n_20753,
       n_20754;
  wire n_20755, n_20756, n_20757, n_20758, n_20759, n_20760, n_20761,
       n_20762;
  wire n_20763, n_20764, n_20765, n_20766, n_20767, n_20768, n_20769,
       n_20770;
  wire n_20771, n_20772, n_20773, n_20774, n_20775, n_20776, n_20777,
       n_20778;
  wire n_20779, n_20780, n_20781, n_20782, n_20783, n_20784, n_20785,
       n_20786;
  wire n_20787, n_20788, n_20789, n_20790, n_20791, n_20792, n_20793,
       n_20794;
  wire n_20795, n_20796, n_20797, n_20798, n_20799, n_20800, n_20801,
       n_20802;
  wire n_20803, n_20804, n_20805, n_20806, n_20807, n_20808, n_20809,
       n_20810;
  wire n_20811, n_20812, n_20813, n_20814, n_20815, n_20816, n_20817,
       n_20818;
  wire n_20819, n_20820, n_20821, n_20822, n_20823, n_20824, n_20825,
       n_20826;
  wire n_20827, n_20828, n_20829, n_20830, n_20831, n_20832, n_20833,
       n_20834;
  wire n_20835, n_20836, n_20837, n_20838, n_20839, n_20840, n_20841,
       n_20842;
  wire n_20843, n_20844, n_20845, n_20846, n_20847, n_20848, n_20849,
       n_20850;
  wire n_20851, n_20852, n_20853, n_20854, n_20855, n_20856, n_20857,
       n_20858;
  wire n_20859, n_20860, n_20861, n_20862, n_20863, n_20864, n_20865,
       n_20866;
  wire n_20867, n_20868, n_20869, n_20870, n_20871, n_20872, n_20873,
       n_20874;
  wire n_20875, n_20876, n_20877, n_20878, n_20879, n_20880, n_20881,
       n_20882;
  wire n_20883, n_20884, n_20885, n_20886, n_20887, n_20888, n_20889,
       n_20890;
  wire n_20891, n_20892, n_20893, n_20894, n_20895, n_20896, n_20897,
       n_20898;
  wire n_20899, n_20900, n_20901, n_20902, n_20903, n_20904, n_20905,
       n_20906;
  wire n_20907, n_20908, n_20909, n_20910;
  CDN_flop \data_stack_mem_reg[0][0] (.clk (clk), .d (n_4684), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [0]));
  CDN_flop \data_stack_mem_reg[0][1] (.clk (clk), .d (n_4688), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [1]));
  CDN_flop \data_stack_mem_reg[0][2] (.clk (clk), .d (n_4692), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [2]));
  CDN_flop \data_stack_mem_reg[0][3] (.clk (clk), .d (n_4696), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [3]));
  CDN_flop \data_stack_mem_reg[0][4] (.clk (clk), .d (n_4700), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [4]));
  CDN_flop \data_stack_mem_reg[0][5] (.clk (clk), .d (n_4704), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [5]));
  CDN_flop \data_stack_mem_reg[0][6] (.clk (clk), .d (n_4708), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [6]));
  CDN_flop \data_stack_mem_reg[0][7] (.clk (clk), .d (n_4712), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [7]));
  CDN_flop \data_stack_mem_reg[1][0] (.clk (clk), .d (n_4716), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [0]));
  CDN_flop \data_stack_mem_reg[1][1] (.clk (clk), .d (n_4720), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [1]));
  CDN_flop \data_stack_mem_reg[1][2] (.clk (clk), .d (n_4724), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [2]));
  CDN_flop \data_stack_mem_reg[1][3] (.clk (clk), .d (n_4728), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [3]));
  CDN_flop \data_stack_mem_reg[1][4] (.clk (clk), .d (n_4732), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [4]));
  CDN_flop \data_stack_mem_reg[1][5] (.clk (clk), .d (n_4736), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [5]));
  CDN_flop \data_stack_mem_reg[1][6] (.clk (clk), .d (n_4740), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [6]));
  CDN_flop \data_stack_mem_reg[1][7] (.clk (clk), .d (n_4744), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [7]));
  CDN_flop \data_stack_mem_reg[2][0] (.clk (clk), .d (n_4748), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [0]));
  CDN_flop \data_stack_mem_reg[2][1] (.clk (clk), .d (n_4752), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [1]));
  CDN_flop \data_stack_mem_reg[2][2] (.clk (clk), .d (n_4756), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [2]));
  CDN_flop \data_stack_mem_reg[2][3] (.clk (clk), .d (n_4760), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [3]));
  CDN_flop \data_stack_mem_reg[2][4] (.clk (clk), .d (n_4764), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [4]));
  CDN_flop \data_stack_mem_reg[2][5] (.clk (clk), .d (n_4768), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [5]));
  CDN_flop \data_stack_mem_reg[2][6] (.clk (clk), .d (n_4772), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [6]));
  CDN_flop \data_stack_mem_reg[2][7] (.clk (clk), .d (n_4776), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [7]));
  CDN_flop \data_stack_mem_reg[3][0] (.clk (clk), .d (n_4780), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [0]));
  CDN_flop \data_stack_mem_reg[3][1] (.clk (clk), .d (n_4784), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [1]));
  CDN_flop \data_stack_mem_reg[3][2] (.clk (clk), .d (n_4788), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [2]));
  CDN_flop \data_stack_mem_reg[3][3] (.clk (clk), .d (n_4792), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [3]));
  CDN_flop \data_stack_mem_reg[3][4] (.clk (clk), .d (n_4796), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [4]));
  CDN_flop \data_stack_mem_reg[3][5] (.clk (clk), .d (n_4800), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [5]));
  CDN_flop \data_stack_mem_reg[3][6] (.clk (clk), .d (n_4804), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [6]));
  CDN_flop \data_stack_mem_reg[3][7] (.clk (clk), .d (n_4808), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [7]));
  CDN_flop \data_stack_mem_reg[4][0] (.clk (clk), .d (n_4812), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [0]));
  CDN_flop \data_stack_mem_reg[4][1] (.clk (clk), .d (n_4816), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [1]));
  CDN_flop \data_stack_mem_reg[4][2] (.clk (clk), .d (n_4820), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [2]));
  CDN_flop \data_stack_mem_reg[4][3] (.clk (clk), .d (n_4824), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [3]));
  CDN_flop \data_stack_mem_reg[4][4] (.clk (clk), .d (n_4828), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [4]));
  CDN_flop \data_stack_mem_reg[4][5] (.clk (clk), .d (n_4832), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [5]));
  CDN_flop \data_stack_mem_reg[4][6] (.clk (clk), .d (n_4836), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [6]));
  CDN_flop \data_stack_mem_reg[4][7] (.clk (clk), .d (n_4840), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [7]));
  CDN_flop \data_stack_mem_reg[5][0] (.clk (clk), .d (n_4844), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [0]));
  CDN_flop \data_stack_mem_reg[5][1] (.clk (clk), .d (n_4848), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [1]));
  CDN_flop \data_stack_mem_reg[5][2] (.clk (clk), .d (n_4852), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [2]));
  CDN_flop \data_stack_mem_reg[5][3] (.clk (clk), .d (n_4856), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [3]));
  CDN_flop \data_stack_mem_reg[5][4] (.clk (clk), .d (n_4860), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [4]));
  CDN_flop \data_stack_mem_reg[5][5] (.clk (clk), .d (n_4864), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [5]));
  CDN_flop \data_stack_mem_reg[5][6] (.clk (clk), .d (n_4868), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [6]));
  CDN_flop \data_stack_mem_reg[5][7] (.clk (clk), .d (n_4872), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [7]));
  CDN_flop \data_stack_mem_reg[6][0] (.clk (clk), .d (n_4876), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [0]));
  CDN_flop \data_stack_mem_reg[6][1] (.clk (clk), .d (n_4880), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [1]));
  CDN_flop \data_stack_mem_reg[6][2] (.clk (clk), .d (n_4884), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [2]));
  CDN_flop \data_stack_mem_reg[6][3] (.clk (clk), .d (n_4888), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [3]));
  CDN_flop \data_stack_mem_reg[6][4] (.clk (clk), .d (n_4892), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [4]));
  CDN_flop \data_stack_mem_reg[6][5] (.clk (clk), .d (n_4896), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [5]));
  CDN_flop \data_stack_mem_reg[6][6] (.clk (clk), .d (n_4900), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [6]));
  CDN_flop \data_stack_mem_reg[6][7] (.clk (clk), .d (n_4904), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [7]));
  CDN_flop \data_stack_mem_reg[7][0] (.clk (clk), .d (n_4908), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [0]));
  CDN_flop \data_stack_mem_reg[7][1] (.clk (clk), .d (n_4912), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [1]));
  CDN_flop \data_stack_mem_reg[7][2] (.clk (clk), .d (n_4916), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [2]));
  CDN_flop \data_stack_mem_reg[7][3] (.clk (clk), .d (n_4920), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [3]));
  CDN_flop \data_stack_mem_reg[7][4] (.clk (clk), .d (n_4924), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [4]));
  CDN_flop \data_stack_mem_reg[7][5] (.clk (clk), .d (n_4928), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [5]));
  CDN_flop \data_stack_mem_reg[7][6] (.clk (clk), .d (n_4932), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [6]));
  CDN_flop \data_stack_mem_reg[7][7] (.clk (clk), .d (n_4936), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [7]));
  CDN_flop \data_stack_mem_reg[8][0] (.clk (clk), .d (n_4940), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [0]));
  CDN_flop \data_stack_mem_reg[8][1] (.clk (clk), .d (n_4944), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [1]));
  CDN_flop \data_stack_mem_reg[8][2] (.clk (clk), .d (n_4948), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [2]));
  CDN_flop \data_stack_mem_reg[8][3] (.clk (clk), .d (n_4952), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [3]));
  CDN_flop \data_stack_mem_reg[8][4] (.clk (clk), .d (n_4956), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [4]));
  CDN_flop \data_stack_mem_reg[8][5] (.clk (clk), .d (n_4960), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [5]));
  CDN_flop \data_stack_mem_reg[8][6] (.clk (clk), .d (n_4964), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [6]));
  CDN_flop \data_stack_mem_reg[8][7] (.clk (clk), .d (n_4968), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [7]));
  CDN_flop \data_stack_pointer_reg[0] (.clk (clk), .d (n_5004), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[0]));
  CDN_flop \data_stack_pointer_reg[1] (.clk (clk), .d (n_5008), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[1]));
  CDN_flop \data_stack_pointer_reg[2] (.clk (clk), .d (n_5012), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[2]));
  CDN_flop \data_stack_pointer_reg[3] (.clk (clk), .d (n_5016), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[3]));
  CDN_flop dout_valid_reg(.clk (clk), .d (n_5019), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (dout_valid));
  not g129 (n_521, rst_n);
  not g1755 (n_523, enable_n);
  nand g17438 (n_12732, out_fifo_read_pointer[1],
       out_fifo_read_pointer[0]);
  nand g18758 (n_12866, n_3902, \data_stack_mem[2] [7]);
  nand g18880 (n_12898, n_3902, \data_stack_mem[2] [2]);
  or g18963 (n_12921, out_fifo_write_pointer[1],
       out_fifo_write_pointer[0]);
  nand g19011 (n_12933, n_3902, \data_stack_mem[2] [4]);
  or g19566 (n_12854, wc, out_fifo_write_pointer[0]);
  not gc (wc, out_fifo_write_pointer[1]);
  or g19567 (n_12847, out_fifo_write_pointer[1], wc0);
  not gc0 (wc0, out_fifo_write_pointer[0]);
  or g19655 (n_12920, n_20, wc1);
  not gc1 (wc1, \data_stack_mem[4] [7]);
  or g19662 (n_12869, n_20, wc2);
  not gc2 (wc2, \data_stack_mem[4] [2]);
  or g19666 (n_12932, n_20, wc3);
  not gc3 (wc3, \data_stack_mem[4] [4]);
  or g19679 (n_12941, n_20, wc4);
  not gc4 (wc4, \data_stack_mem[4] [1]);
  nand g26004 (n_13400, data_stack_pointer[3], \data_stack_mem[7] [1]);
  nand g26010 (n_13401, data_stack_pointer[3], \data_stack_mem[7] [7]);
  nand g26016 (n_13402, data_stack_pointer[3], \data_stack_mem[7] [2]);
  nand g26022 (n_13403, data_stack_pointer[3], \data_stack_mem[7] [4]);
  nand g27145 (n_12917, n_3902, \data_stack_mem[2] [1]);
  or g27618 (n_13409, n_1425, wc5);
  not gc5 (wc5, \data_stack_mem[8] [0]);
  or g27753 (n_4634, n_3793, data_stack_pointer[0]);
  or g30837 (n_13778, enable_n, sh_bit_cnt[0]);
  nand g30889 (n_13789, data_stack_pointer[1], data_stack_pointer[0]);
  or g30897 (n_13215, out_fifo_write_pointer[2], n_131);
  or g30928 (n_13214, wc6, n_131);
  not gc6 (wc6, out_fifo_write_pointer[2]);
  nand g30936 (n_13798, n_1361, \data_stack_mem[4] [0]);
  nand g30948 (n_13803, n_3902, \data_stack_mem[2] [3]);
  nand g30957 (n_13805, n_1377, \data_stack_mem[5] [0]);
  or g30961 (n_13806, sh_bit_cnt[1], n_13778);
  nand g30969 (n_13807, n_1393, \data_stack_mem[6] [0]);
  nand g30995 (n_13811, n_1329, \data_stack_mem[2] [0]);
  nand g30999 (n_13812, n_1345, \data_stack_mem[3] [0]);
  nand g31003 (n_13813, n_1409, \data_stack_mem[7] [0]);
  or g31012 (n_13815, sh_reg_out_bit_counter[1],
       sh_reg_out_bit_counter[0]);
  or g31066 (n_13827, wc7, n_13203);
  not gc7 (wc7, n_4209);
  or g31332 (n_13906, n_12809, n_4369);
  nand g31338 (n_170, n_13907, n_13792);
  nand g31354 (n_13912, n_3902, \data_stack_mem[2] [5]);
  nand g31371 (n_13916, \data_stack_mem[1] [0], \data_stack_mem[0] [0]);
  nand g31378 (n_13918, \data_stack_mem[1] [4], \data_stack_mem[0] [4]);
  nand g31382 (n_13919, \data_stack_mem[1] [2], \data_stack_mem[0] [2]);
  nand g31388 (n_13428, n_13920, n_13795);
  nand g31390 (n_13921, n_1425, \data_stack_mem[8] [0]);
  or g31434 (n_13932, data_stack_pointer[2], data_stack_pointer[1]);
  or g31438 (n_13933, sh_reg_in[1], sh_reg_in[0]);
  or g31442 (n_13934, sh_reg_out_bit_counter[2], n_13815);
  or g31443 (n_13121, n_13934, sh_reg_out_bit_counter[3]);
  nand g31448 (n_1326, n_13935, n_13780);
  or g31450 (n_13936, n_13141, n_4433);
  or g31451 (n_12905, n_13936, n_4432);
  nand g31459 (n_13938, \data_stack_mem[1] [6], \data_stack_mem[0] [6]);
  or g31488 (n_13439, n_13945, n_13147);
  or g31490 (n_13946, n_12921, n_13214);
  not g31492 (n_847, n_13946);
  or g31494 (n_13947, n_12854, n_13214);
  not g31496 (n_827, n_13947);
  or g31498 (n_13948, data_stack_pointer[3], data_stack_pointer[1]);
  or g31502 (n_13949, n_12847, n_13215);
  not g31504 (n_877, n_13949);
  or g31510 (n_13951, n_12854, n_13215);
  not g31512 (n_867, n_13951);
  or g31529 (n_13956, n_12847, n_13214);
  not g31531 (n_837, n_13956);
  nand g31536 (n_13958, data_stack_pointer[3], \data_stack_mem[7] [5]);
  nand g31540 (n_13959, data_stack_pointer[3], \data_stack_mem[7] [6]);
  or g31544 (n_13960, n_13146, n_4497);
  or g31545 (n_12860, n_13960, n_4496);
  or g31548 (n_13961, n_12921, n_13215);
  not g31550 (n_887, n_13961);
  or g31558 (n_13964, wc8, n_20);
  not gc8 (wc8, \data_stack_mem[4] [3]);
  nand g31562 (n_13965, data_stack_pointer[3], \data_stack_mem[7] [3]);
  or g31589 (n_13972, n_12814, n_4401);
  nand g31611 (n_13978, n_3902, \data_stack_mem[2] [6]);
  or g32176 (n_13814, wc9, \data_stack_mem[0] [0]);
  not gc9 (wc9, \data_stack_mem[1] [0]);
  or g32178 (n_13907, \data_stack_mem[1] [2], wc10);
  not gc10 (wc10, \data_stack_mem[0] [2]);
  or g32181 (n_13920, \data_stack_mem[1] [4], wc11);
  not gc11 (wc11, \data_stack_mem[0] [4]);
  or g32184 (n_13935, wc12, \data_stack_mem[0] [6]);
  not gc12 (wc12, \data_stack_mem[1] [6]);
  or g32189 (n_13903, data_stack_pointer[3], wc13);
  not gc13 (wc13, data_stack_pointer[0]);
  or g32190 (n_13942, data_stack_pointer[3], wc14);
  not gc14 (wc14, data_stack_pointer[2]);
  or g32216 (n_13825, wc15, \data_stack_mem[2] [1]);
  not gc15 (wc15, n_3902);
  or g32223 (n_13821, wc16, \data_stack_mem[2] [5]);
  not gc16 (wc16, n_3902);
  or g32234 (n_13966, n_20, wc17);
  not gc17 (wc17, \data_stack_mem[4] [5]);
  or g32238 (n_13970, n_20, wc18);
  not gc18 (wc18, \data_stack_mem[4] [6]);
  or g32271 (n_131, n_158, wc19);
  not gc19 (wc19, sh_reg_in[8]);
  or g32276 (n_13784, n_1329, wc20);
  not gc20 (wc20, \data_stack_mem[2] [0]);
  or g32323 (n_13788, n_1345, wc21);
  not gc21 (wc21, \data_stack_mem[3] [0]);
  or g32399 (n_13779, n_1361, wc22);
  not gc22 (wc22, \data_stack_mem[4] [0]);
  or g32433 (n_13781, n_1377, wc23);
  not gc23 (wc23, \data_stack_mem[5] [0]);
  or g32447 (n_13783, n_1393, wc24);
  not gc24 (wc24, \data_stack_mem[6] [0]);
  or g32463 (n_13791, n_1409, wc25);
  not gc25 (wc25, \data_stack_mem[7] [0]);
  or g32490 (n_14063, n_12824, wc26);
  not gc26 (wc26, n_4081);
  or g32511 (n_13809, n_12813, wc27);
  not gc27 (wc27, n_4113);
  or g32531 (n_13822, n_13220, wc28);
  not gc28 (wc28, n_4145);
  or g32547 (n_13914, n_13197, wc29);
  not gc29 (wc29, n_4177);
  or g32576 (n_13931, n_13439, wc30);
  not gc30 (wc30, n_4240);
  or g33469 (n_14171, \data_stack_mem[1] [3], \data_stack_mem[0] [3]);
  or g33472 (n_14172, \data_stack_mem[1] [5], \data_stack_mem[0] [5]);
  or g33488 (n_14178, n_13121, sh_reg_out_bit_counter[4]);
  or g33501 (n_13794, \data_stack_mem[1] [4], \data_stack_mem[0] [4]);
  or g33504 (n_14184, n_13933, sh_reg_in[4]);
  or g33510 (n_13774, \data_stack_mem[1] [6], \data_stack_mem[0] [6]);
  or g33513 (n_13793, \data_stack_mem[1] [2], \data_stack_mem[0] [2]);
  or g33537 (n_14195, n_11641, \data_stack_mem[5] [4]);
  or g33543 (n_14197, n_11576, \data_stack_mem[4] [5]);
  or g33546 (n_14198, wc31, n_12170);
  not gc31 (wc31, \data_stack_mem[4] [5]);
  or g33552 (n_14200, wc32, n_13783);
  not gc32 (wc32, \data_stack_mem[6] [1]);
  or g33555 (n_14201, wc33, n_12265);
  not gc33 (wc33, \data_stack_mem[5] [3]);
  or g33558 (n_14202, n_11673, \data_stack_mem[5] [3]);
  or g33561 (n_14203, wc34, n_12076);
  not gc34 (wc34, \data_stack_mem[3] [6]);
  or g33564 (n_14204, n_11480, \data_stack_mem[3] [6]);
  or g33567 (n_14205, n_11540, \data_stack_mem[4] [4]);
  or g33570 (n_14206, n_11622, \data_stack_mem[5] [2]);
  or g33573 (n_14207, wc35, n_12141);
  not gc35 (wc35, \data_stack_mem[4] [4]);
  or g33576 (n_14208, wc36, n_12218);
  not gc36 (wc36, \data_stack_mem[5] [2]);
  or g33582 (n_14210, wc37, n_12725);
  not gc37 (wc37, \data_stack_mem[2] [7]);
  nand g33585 (n_14211, n_12648, \data_stack_mem[2] [7]);
  or g33588 (n_14212, n_11572, \data_stack_mem[4] [3]);
  or g33591 (n_14213, n_11478, \data_stack_mem[3] [5]);
  or g33594 (n_14214, wc38, n_12074);
  not gc38 (wc38, \data_stack_mem[3] [5]);
  or g33600 (n_14216, wc39, n_13781);
  not gc39 (wc39, \data_stack_mem[5] [1]);
  or g33603 (n_14217, wc40, n_12166);
  not gc40 (wc40, \data_stack_mem[4] [3]);
  or g33612 (n_14220, n_11521, \data_stack_mem[4] [2]);
  or g33615 (n_14221, \data_stack_mem[3] [4], n_11449);
  or g33618 (n_14222, wc41, n_12045);
  not gc41 (wc41, \data_stack_mem[3] [4]);
  or g33621 (n_14223, wc42, n_12119);
  not gc42 (wc42, \data_stack_mem[4] [2]);
  or g33624 (n_14224, n_12645, \data_stack_mem[2] [6]);
  or g33627 (n_14225, wc43, n_12722);
  not gc43 (wc43, \data_stack_mem[2] [6]);
  or g33633 (n_14227, wc44, n_12070);
  not gc44 (wc44, \data_stack_mem[3] [3]);
  or g33639 (n_14229, n_11980, \data_stack_mem[8] [5]);
  or g33642 (n_14230, wc45, n_12240);
  not gc45 (wc45, \data_stack_mem[5] [4]);
  or g33645 (n_14231, n_12643, \data_stack_mem[2] [5]);
  or g33648 (n_14232, \data_stack_mem[2] [1], wc46);
  not gc46 (wc46, n_13811);
  or g33651 (n_14233, n_11723, \data_stack_mem[6] [2]);
  or g33654 (n_14234, \data_stack_mem[3] [2], n_11432);
  or g33659 (n_14236, wc47, n_12317);
  not gc47 (wc47, \data_stack_mem[6] [2]);
  or g33665 (n_14238, n_11578, \data_stack_mem[4] [6]);
  or g33674 (n_14242, n_13788, n_4376);
  or g33680 (n_14244, wc48, n_12683);
  not gc48 (wc48, \data_stack_mem[2] [2]);
  nand g33685 (n_14246, n_3902, \data_stack_mem[2] [0]);
  or g33688 (n_14247, wc49, n_12172);
  not gc49 (wc49, \data_stack_mem[4] [6]);
  nand g33691 (n_14248, \data_stack_mem[3] [7], n_11483);
  or g33694 (n_14249, wc50, n_12699);
  not gc50 (wc50, \data_stack_mem[2] [4]);
  or g33697 (n_14250, wc51, n_12467);
  not gc51 (wc51, \data_stack_mem[7] [5]);
  or g33702 (n_14252, n_11881, \data_stack_mem[7] [6]);
  nand g33705 (n_14253, n_11783, \data_stack_mem[6] [7]);
  or g33707 (n_14060, wc52, n_14228);
  not gc52 (wc52, n_14253);
  or g33708 (n_14254, wc53, n_12373);
  not gc53 (wc53, \data_stack_mem[6] [7]);
  or g33711 (n_14255, wc54, n_12469);
  not gc54 (wc54, \data_stack_mem[7] [6]);
  or g33714 (n_14256, wc55, n_12269);
  not gc55 (wc55, \data_stack_mem[5] [5]);
  or g33720 (n_14258, n_12622, \data_stack_mem[2] [4]);
  or g33723 (n_14259, wc56, n_4534);
  not gc56 (wc56, \data_stack_mem[8] [3]);
  or g33726 (n_14260, wc57, n_12416);
  not gc57 (wc57, \data_stack_mem[7] [2]);
  or g33729 (n_14261, n_11879, \data_stack_mem[7] [5]);
  or g33732 (n_14262, n_4245, \data_stack_mem[8] [4]);
  or g33738 (n_14264, n_11982, \data_stack_mem[8] [6]);
  or g33741 (n_14265, wc58, n_13791);
  not gc58 (wc58, \data_stack_mem[7] [1]);
  or g33744 (n_14266, n_13784, n_4344);
  or g33747 (n_14267, n_13827, wc59);
  not gc59 (wc59, n_4208);
  or g33750 (n_14268, wc60, n_12339);
  not gc60 (wc60, \data_stack_mem[6] [4]);
  or g33753 (n_14269, n_4054, n_12639);
  or g33756 (n_14270, wc61, n_13779);
  not gc61 (wc61, \data_stack_mem[4] [1]);
  or g33759 (n_14271, wc62, n_4532);
  not gc62 (wc62, \data_stack_mem[8] [5]);
  or g33762 (n_14272, wc63, n_4531);
  not gc63 (wc63, \data_stack_mem[8] [6]);
  or g33765 (n_14273, wc64, n_12720);
  not gc64 (wc64, \data_stack_mem[2] [5]);
  or g33768 (n_14274, wc65, n_12175);
  not gc65 (wc65, \data_stack_mem[4] [7]);
  nand g33771 (n_14275, n_11884, \data_stack_mem[7] [7]);
  or g33774 (n_14276, n_11824, \data_stack_mem[7] [2]);
  nand g33777 (n_14277, n_4242, \data_stack_mem[8] [7]);
  or g33780 (n_14278, wc66, n_12472);
  not gc66 (wc66, \data_stack_mem[7] [7]);
  nand g33783 (n_14279, n_11682, \data_stack_mem[5] [7]);
  or g33789 (n_14281, n_13806, sh_bit_cnt[2]);
  or g33790 (n_158, n_14281, sh_bit_cnt[3]);
  or g33792 (n_14282, n_11875, \data_stack_mem[7] [3]);
  or g33795 (n_14283, n_4501, n_12438);
  or g33798 (n_14284, wc67, n_12716);
  not gc67 (wc67, \data_stack_mem[2] [3]);
  or g33806 (n_14287, n_11976, \data_stack_mem[8] [3]);
  or g33809 (n_14288, n_4375, n_12027);
  or g33812 (n_14289, n_12606, \data_stack_mem[2] [2]);
  or g33815 (n_14290, n_11774, \data_stack_mem[6] [3]);
  or g33818 (n_14291, wc68, n_4216);
  not gc68 (wc68, n_13813);
  or g33821 (n_14292, n_11474, \data_stack_mem[3] [3]);
  or g33824 (n_14293, wc69, n_12364);
  not gc69 (wc69, \data_stack_mem[6] [3]);
  nand g33827 (n_14294, n_3793, \data_stack_mem[1] [0]);
  or g33836 (n_14297, \data_stack_mem[1] [1], \data_stack_mem[0] [1]);
  or g33839 (n_14298, n_4247, \data_stack_mem[8] [2]);
  or g33842 (n_14299, n_11679, \data_stack_mem[5] [6]);
  or g33854 (n_14303, n_4248, \data_stack_mem[8] [1]);
  or g33857 (n_14304, wc70, n_12370);
  not gc70 (wc70, \data_stack_mem[6] [6]);
  or g33860 (n_14305, wc71, n_12274);
  not gc71 (wc71, \data_stack_mem[5] [7]);
  or g33862 (n_14045, wc72, n_14280);
  not gc72 (wc72, n_14305);
  or g33865 (n_14307, n_11843, \data_stack_mem[7] [4]);
  or g33868 (n_14308, wc73, n_12463);
  not gc73 (wc73, \data_stack_mem[7] [3]);
  or g33871 (n_14309, n_11780, \data_stack_mem[6] [6]);
  or g33874 (n_14310, n_11778, \data_stack_mem[6] [5]);
  or g33877 (n_14311, n_11677, \data_stack_mem[5] [5]);
  or g33880 (n_14312, n_11742, \data_stack_mem[6] [4]);
  or g33883 (n_14313, wc74, n_12271);
  not gc74 (wc74, \data_stack_mem[5] [6]);
  or g33886 (n_14314, wc75, n_12368);
  not gc75 (wc75, \data_stack_mem[6] [5]);
  or g33889 (n_14315, wc76, n_12079);
  not gc76 (wc76, \data_stack_mem[3] [7]);
  nand g33892 (n_14316, n_11581, \data_stack_mem[4] [7]);
  or g33894 (n_14085, wc77, n_14286);
  not gc77 (wc77, n_14316);
  or g33898 (n_14296, wc78, \data_stack_mem[0] [1]);
  not gc78 (wc78, \data_stack_mem[1] [1]);
  or g33899 (n_13792, wc79, \data_stack_mem[0] [2]);
  not gc79 (wc79, \data_stack_mem[1] [2]);
  or g33900 (n_14175, wc80, \data_stack_mem[0] [3]);
  not gc80 (wc80, \data_stack_mem[1] [3]);
  or g33901 (n_13795, wc81, \data_stack_mem[0] [4]);
  not gc81 (wc81, \data_stack_mem[1] [4]);
  or g33902 (n_14174, wc82, \data_stack_mem[0] [5]);
  not gc82 (wc82, \data_stack_mem[1] [5]);
  or g33903 (n_13780, \data_stack_mem[1] [6], wc83);
  not gc83 (wc83, \data_stack_mem[0] [6]);
  or g33904 (n_14170, \data_stack_mem[1] [7], wc84);
  not gc84 (wc84, \data_stack_mem[0] [7]);
  or g33914 (n_14226, n_20, wc85);
  not gc85 (wc85, \data_stack_mem[4] [0]);
  or g33917 (n_14302, n_11331, wc86);
  not gc86 (wc86, \data_stack_mem[8] [0]);
  or g33951 (n_14243, wc87, \data_stack_mem[3] [1]);
  not gc87 (wc87, n_13812);
  or g33984 (n_14263, wc88, \data_stack_mem[4] [1]);
  not gc88 (wc88, n_13798);
  or g33998 (n_14215, wc89, \data_stack_mem[5] [1]);
  not gc89 (wc89, n_13805);
  or g34016 (n_14199, wc90, \data_stack_mem[6] [1]);
  not gc90 (wc90, n_13807);
  or g34064 (n_14116, n_14218, wc91);
  not gc91 (wc91, n_14210);
  or g34078 (n_14075, n_14219, wc92);
  not gc92 (wc92, n_14211);
  or g34130 (n_14038, n_14317, wc93);
  not gc93 (wc93, n_14274);
  or g34147 (n_14030, n_14300, wc94);
  not gc94 (wc94, n_14279);
  or g34150 (n_14257, n_13809, wc95);
  not gc95 (wc95, n_4112);
  or g34165 (n_14181, n_13822, wc96);
  not gc96 (wc96, n_4144);
  or g34169 (n_14058, n_14295, wc97);
  not gc97 (wc97, n_14254);
  or g34176 (n_14301, n_13914, wc98);
  not gc98 (wc98, n_4176);
  or g34243 (n_13928, n_12895, wc99);
  not gc99 (wc99, n_4049);
  nand g34448 (n_14470, n_13131, n_14191);
  or g34451 (n_14471, wc100, n_12571);
  not gc100 (wc100, \data_stack_mem[8] [7]);
  nand g34469 (n_14480, n_13443, n_14190);
  or g34512 (n_14501, wc101, n_4533);
  not gc101 (wc101, \data_stack_mem[8] [4]);
  nand g34542 (n_14516, n_3793, n_13794);
  or g34552 (n_14521, wc102, n_12515);
  not gc102 (wc102, \data_stack_mem[8] [2]);
  nand g34558 (n_14524, \data_stack_mem[7] [0], data_stack_pointer[3]);
  or g34564 (n_14527, n_13409, wc103);
  not gc103 (wc103, \data_stack_mem[8] [1]);
  nand g34582 (n_14536, n_3793, n_13793);
  or g34600 (n_14545, wc104, data_stack_pointer[3]);
  not gc104 (wc104, n_13789);
  nand g34610 (n_14550, n_3793, n_14297);
  or g34622 (n_14556, n_13903, wc105);
  not gc105 (wc105, data_stack_pointer[2]);
  or g34626 (n_14558, wc106, data_stack_pointer[2]);
  not gc106 (wc106, data_stack_pointer[0]);
  or g34660 (n_14575, \data_stack_mem[8] [0], n_11331);
  or g34678 (n_14584, n_100, n_12732);
  or g34721 (n_14566, n_14621, n_14622);
  or g38691 (n_14191, wc107, result[8]);
  not gc107 (wc107, result[12]);
  or g38693 (n_14190, wc108, result[9]);
  not gc108 (wc108, result[12]);
  nand g38695 (n_5763, n_19298, n_19299);
  nand g38696 (n_5771, n_19304, n_19305);
  nand g38697 (n_5747, n_19310, n_19311);
  nand g38698 (n_5775, n_19340, n_19341);
  nand g38699 (n_5767, n_19322, n_19323);
  nand g38700 (n_5759, n_19328, n_19329);
  nand g38701 (n_5755, n_19334, n_19335);
  nand g38702 (n_5751, n_19316, n_19317);
  or g38703 (n_19340, wc109, n_12775);
  not gc109 (wc109, n_633);
  or g38704 (n_19304, wc110, n_12766);
  not gc110 (wc110, n_633);
  or g38705 (n_19322, wc111, n_12769);
  not gc111 (wc111, n_633);
  or g38706 (n_19334, wc112, n_12774);
  not gc112 (wc112, n_633);
  or g38707 (n_19298, wc113, n_12765);
  not gc113 (wc113, n_633);
  or g38708 (n_19310, wc114, n_12767);
  not gc114 (wc114, n_633);
  or g38709 (n_19328, wc115, n_12772);
  not gc115 (wc115, n_633);
  or g38710 (n_19316, wc116, n_12768);
  not gc116 (wc116, n_633);
  nand g38711 (n_5719, n_19268, n_19269);
  nand g38712 (n_5723, n_19286, n_19287);
  nand g38713 (n_5731, n_19250, n_19251);
  or g38714 (n_20604, wc117, n_4646);
  not gc117 (wc117, n_4643);
  or g38715 (n_20605, n_4643, wc118);
  not gc118 (wc118, n_4646);
  nand g38716 (n_633, n_20604, n_20605);
  nand g38717 (n_5739, n_19256, n_19257);
  nand g38718 (n_5727, n_19280, n_19281);
  nand g38719 (n_5715, n_19262, n_19263);
  nand g38720 (n_5735, n_19274, n_19275);
  nand g38721 (n_5743, n_19292, n_19293);
  or g38722 (n_19292, wc119, n_12775);
  not gc119 (wc119, n_624);
  or g38723 (n_19280, wc120, n_12772);
  not gc120 (wc120, n_624);
  or g38724 (n_19268, wc121, n_12768);
  not gc121 (wc121, n_624);
  or g38725 (n_20606, wc122, n_4642);
  not gc122 (wc122, n_14470);
  or g38726 (n_20607, n_14470, wc123);
  not gc123 (wc123, n_4642);
  nand g38727 (n_4643, n_20606, n_20607);
  or g38728 (n_19250, wc124, n_12765);
  not gc124 (wc124, n_624);
  or g38729 (n_19286, wc125, n_12774);
  not gc125 (wc125, n_624);
  or g38730 (n_19262, wc126, n_12767);
  not gc126 (wc126, n_624);
  or g38731 (n_19256, wc127, n_12766);
  not gc127 (wc127, n_624);
  or g38732 (n_19274, wc128, n_12769);
  not gc128 (wc128, n_624);
  nand g38733 (n_5495, n_19130, n_19131);
  nand g38734 (n_5567, n_19166, n_19167);
  nand g38735 (n_4642, n_19244, n_19245);
  nand g38736 (n_5435, n_19106, n_19107);
  nand g38737 (n_5291, n_19232, n_19233);
  nand g38738 (n_5135, n_19142, n_19143);
  nand g38739 (n_5279, n_19154, n_19155);
  nand g38740 (n_5063, n_19136, n_19137);
  nand g38741 (n_5147, n_19094, n_19095);
  nand g38742 (n_5507, n_19070, n_19071);
  nand g38743 (n_5579, n_19238, n_19239);
  or g38744 (n_20608, wc129, n_4640);
  not gc129 (wc129, n_4637);
  or g38745 (n_20609, n_4637, wc130);
  not gc130 (wc130, n_4640);
  nand g38746 (n_624, n_20608, n_20609);
  nand g38747 (n_5351, n_19124, n_19125);
  nand g38748 (n_5363, n_19058, n_19059);
  nand g38749 (n_5075, n_19082, n_19083);
  nand g38753 (n_5207, n_19160, n_19161);
  nand g38754 (n_5423, n_19148, n_19149);
  nand g38755 (n_5219, n_19118, n_19119);
  or g38756 (n_19166, n_12775, wc131);
  not gc131 (wc131, result[7]);
  or g38757 (n_19136, n_12767, wc132);
  not gc132 (wc132, result[7]);
  or g38758 (n_19238, n_12775, wc133);
  not gc133 (wc133, result[10]);
  or g38759 (n_19058, n_12765, wc134);
  not gc134 (wc134, result[10]);
  nand g38760 (n_5503, n_19064, n_19065);
  or g38761 (n_19232, n_12772, wc135);
  not gc135 (wc135, result[10]);
  nand g38762 (n_5575, n_19226, n_19227);
  nand g38763 (n_5359, n_19052, n_19053);
  or g38764 (n_19160, n_12774, wc136);
  not gc136 (wc136, result[7]);
  nand g38765 (n_5287, n_19220, n_19221);
  or g38766 (n_19070, n_12766, wc137);
  not gc137 (wc137, result[10]);
  or g38767 (n_19130, n_12766, wc138);
  not gc138 (wc138, result[7]);
  or g38768 (n_19244, wc139, result[10]);
  not gc139 (wc139, result[12]);
  or g38769 (n_19142, n_12768, wc140);
  not gc140 (wc140, result[7]);
  or g38770 (n_19124, n_12765, wc141);
  not gc141 (wc141, result[7]);
  nand g38771 (n_5071, n_19076, n_19077);
  or g38772 (n_19082, n_12767, wc142);
  not gc142 (wc142, result[10]);
  or g38773 (n_19154, n_12772, wc143);
  not gc143 (wc143, result[7]);
  or g38774 (n_19118, n_12774, wc144);
  not gc144 (wc144, result[10]);
  nand g38775 (n_5215, n_19112, n_19113);
  nand g38776 (n_5143, n_19088, n_19089);
  or g38777 (n_19094, n_12768, wc145);
  not gc145 (wc145, result[10]);
  or g38778 (n_20612, wc146, result[7]);
  not gc146 (wc146, n_13909);
  or g38779 (n_20613, n_13909, wc147);
  not gc147 (wc147, result[7]);
  nand g38780 (n_4637, n_20612, n_20613);
  or g38781 (n_19148, n_12769, wc148);
  not gc148 (wc148, result[7]);
  nand g38782 (n_5431, n_19100, n_19101);
  or g38783 (n_19106, n_12769, wc149);
  not gc149 (wc149, result[10]);
  or g38784 (n_19112, n_12774, wc150);
  not gc150 (wc150, result[9]);
  or g38785 (n_19100, n_12769, wc151);
  not gc151 (wc151, result[9]);
  or g38786 (n_19088, n_12768, wc152);
  not gc152 (wc152, result[9]);
  nand g38787 (n_5211, n_18902, n_18903);
  nand g38788 (n_5427, n_18896, n_18897);
  or g38789 (n_19076, n_12767, wc153);
  not gc153 (wc153, result[9]);
  nand g38790 (n_5139, n_18890, n_18891);
  or g38791 (n_19220, wc154, n_12772);
  not gc154 (wc154, result[9]);
  or g38792 (n_19226, wc155, n_12775);
  not gc155 (wc155, result[9]);
  nand g38793 (n_5067, n_18884, n_18885);
  nand g38794 (n_5499, n_18878, n_18879);
  or g38795 (n_19064, n_12766, wc156);
  not gc156 (wc156, result[9]);
  nand g38796 (n_5355, n_18872, n_18873);
  or g38797 (result[10], wc157, n_19611);
  not gc157 (wc157, n_19245);
  or g38798 (n_19052, n_12765, wc158);
  not gc158 (wc158, result[9]);
  nand g38799 (n_5571, n_19010, n_19011);
  or g38800 (result[7], n_19046, n_19047);
  nand g38801 (n_5283, n_19004, n_19005);
  nand g38802 (n_5371, n_13988, n_18951);
  nand g38803 (n_5379, n_13988, n_18948);
  nand g38804 (n_5375, n_13988, n_18945);
  nand g38805 (n_5095, n_13990, n_18954);
  nand g38806 (n_5383, n_13988, n_18942);
  nand g38807 (n_5447, n_13985, n_18939);
  nand g38808 (n_5087, n_13990, n_18957);
  nand g38809 (n_5451, n_13985, n_18936);
  nand g38810 (n_5455, n_13985, n_18933);
  nand g38811 (n_5091, n_13990, n_18960);
  nand g38812 (n_5583, n_19172, n_19173);
  nand g38813 (n_5443, n_13985, n_18930);
  nand g38814 (n_5083, n_13990, n_18963);
  nand g38815 (n_5595, n_13984, n_18927);
  nand g38816 (n_5223, n_19178, n_19179);
  nand g38817 (n_5163, n_13991, n_18966);
  nand g38818 (n_5591, n_13984, n_18924);
  nand g38819 (n_5587, n_13984, n_18921);
  nand g38820 (n_5155, n_13991, n_18969);
  nand g38821 (n_5295, n_19184, n_19185);
  nand g38822 (n_5599, n_13984, n_18918);
  nand g38823 (n_5167, n_13991, n_18972);
  nand g38824 (n_5515, n_13983, n_18915);
  or g38825 (n_19004, n_12772, wc159);
  not gc159 (wc159, result[8]);
  nand g38826 (n_5159, n_13991, n_18975);
  nand g38827 (n_5519, n_13983, n_18912);
  nand g38828 (n_5527, n_13983, n_18909);
  nand g38829 (n_5311, n_13993, n_18978);
  nand g38830 (n_5151, n_19196, n_19197);
  nand g38831 (n_5523, n_13983, n_18906);
  nand g38832 (n_5299, n_13993, n_18981);
  nand g38833 (n_5079, n_19202, n_19203);
  or g38834 (n_18902, n_12774, wc160);
  not gc160 (wc160, result[8]);
  nand g38835 (n_5303, n_13993, n_18984);
  nand g38836 (n_5511, n_19208, n_19209);
  or g38837 (n_18896, n_12769, wc161);
  not gc161 (wc161, result[8]);
  nand g38838 (n_5307, n_13993, n_18987);
  nand g38839 (n_5367, n_19214, n_19215);
  or g38840 (n_18890, n_12768, wc162);
  not gc162 (wc162, result[8]);
  nand g38841 (n_5235, n_13994, n_18990);
  or g38842 (n_18884, n_12767, wc163);
  not gc163 (wc163, result[8]);
  or g38843 (n_18878, n_12766, wc164);
  not gc164 (wc164, result[8]);
  nand g38844 (n_5231, n_13994, n_18993);
  or g38845 (n_18872, n_12765, wc165);
  not gc165 (wc165, result[8]);
  nand g38846 (n_5239, n_13994, n_18996);
  nand g38847 (n_19611, n_19609, n_19610);
  or g38848 (result[9], n_19020, wc166);
  not gc166 (wc166, n_13443);
  nand g38849 (n_5227, n_13994, n_18999);
  or g38850 (n_19010, n_12775, wc167);
  not gc167 (wc167, result[8]);
  nand g38851 (n_19046, n_19042, n_19043);
  nand g38852 (n_5439, n_19190, n_19191);
  nand g38853 (n_5347, n_18791, n_18792);
  or g38854 (n_13985, n_12847, n_13777);
  or g38855 (n_19196, wc168, n_12768);
  not gc168 (wc168, n_13775);
  nand g38856 (n_5203, n_18827, n_18828);
  or g38857 (result[8], wc169, n_18867);
  not gc169 (wc169, n_14141);
  or g38858 (n_13988, n_12921, n_13777);
  or g38859 (n_19202, wc170, n_12767);
  not gc170 (wc170, n_13775);
  nand g38860 (n_5275, n_18821, n_18822);
  nand g38861 (n_20614, n_13915, n_13772);
  or g38862 (n_20615, n_13915, n_13772);
  nand g38863 (n_4640, n_20614, n_20615);
  or g38864 (n_19208, wc171, n_12766);
  not gc171 (wc171, n_13775);
  or g38865 (n_13993, n_139, n_13776);
  nand g38866 (n_5419, n_18815, n_18816);
  or g38867 (n_19214, wc172, n_12765);
  not gc172 (wc172, n_13775);
  or g38868 (n_13994, n_12854, n_13776);
  or g38869 (n_13990, n_12921, n_13776);
  or g38870 (n_19172, wc173, n_12775);
  not gc173 (wc173, n_13775);
  nand g38871 (n_5131, n_18809, n_18810);
  nand g38872 (n_19042, n_4634, n_3676);
  nand g38873 (n_19020, n_19018, n_19019);
  or g38874 (n_19178, wc174, n_12774);
  not gc174 (wc174, n_13775);
  nand g38875 (n_5059, n_18803, n_18804);
  or g38876 (n_13991, n_12847, n_13776);
  nand g38877 (n_19610, n_13782, n_14472);
  or g38878 (n_19184, wc175, n_12772);
  not gc175 (wc175, n_13775);
  nand g38879 (n_5491, n_18797, n_18798);
  or g38880 (n_13983, n_12854, n_13777);
  or g38881 (n_13984, n_139, n_13777);
  or g38882 (n_19190, wc176, n_12769);
  not gc176 (wc176, n_13775);
  nand g38883 (n_5563, n_18833, n_18834);
  or g38884 (n_18815, n_12769, wc177);
  not gc177 (wc177, result[6]);
  or g38885 (n_14472, n_12853, wc178);
  not gc178 (wc178, n_18852);
  or g38886 (n_13777, n_18846, wc179);
  not gc179 (wc179, rst_n);
  or g38887 (n_18821, n_12772, wc180);
  not gc180 (wc180, result[6]);
  or g38888 (n_13775, result[12], wc181);
  not gc181 (wc181, n_3649);
  nand g38889 (n_20616, result[6], result[1]);
  or g38890 (n_20617, result[6], result[1]);
  nand g38891 (n_13772, n_20616, n_20617);
  or g38892 (n_18827, n_12774, wc182);
  not gc182 (wc182, result[6]);
  nand g38893 (n_18867, n_13131, n_18866);
  or g38894 (n_18833, n_12775, wc183);
  not gc183 (wc183, result[6]);
  nand g38895 (n_19019, n_4528, n_12853);
  or g38896 (n_18791, n_12765, wc184);
  not gc184 (wc184, result[6]);
  or g38897 (n_18797, n_12766, wc185);
  not gc185 (wc185, result[6]);
  or g38898 (n_18803, n_12767, wc186);
  not gc186 (wc186, result[6]);
  or g38899 (n_3676, wc187, n_13190);
  not gc187 (wc187, n_14465);
  or g38900 (n_13776, n_18849, wc188);
  not gc188 (wc188, rst_n);
  or g38901 (n_19609, n_13782, n_19018);
  or g38902 (n_18809, n_12768, wc189);
  not gc189 (wc189, result[6]);
  nand g38903 (n_18866, n_4529, n_14189);
  or g38904 (n_18849, n_13215, wc190);
  not gc190 (wc190, result[12]);
  or g38905 (n_18846, n_13214, wc191);
  not gc191 (wc191, result[12]);
  or g38906 (n_19018, n_4528, n_14141);
  or g38907 (n_12853, n_14189, wc192);
  not gc192 (wc192, n_18843);
  or g38908 (result[6], n_18785, n_18786);
  or g38909 (n_19245, wc193, n_3634);
  not gc193 (wc193, n_2033);
  or g38910 (n_13443, n_18858, n_3634);
  or g38911 (n_13190, wc194, n_3669);
  not gc194 (wc194, n_14464);
  or g38912 (n_3649, n_18861, n_3634);
  nand g38913 (n_5559, n_18722, n_18723);
  nand g38914 (n_3669, n_18746, n_18747);
  or g38915 (n_13131, n_18840, n_3634);
  nand g38916 (n_5199, n_18716, n_18717);
  or g38917 (n_18786, wc195, n_18784);
  not gc195 (wc195, n_18783);
  nand g38918 (n_5271, n_18710, n_18711);
  nand g38919 (n_5415, n_18704, n_18705);
  nand g38920 (n_5127, n_18698, n_18699);
  nand g38921 (n_5055, n_18692, n_18693);
  nand g38922 (n_5487, n_18686, n_18687);
  nand g38923 (n_5343, n_18680, n_18681);
  nand g38924 (result[12], n_18758, n_18759);
  or g38925 (n_14141, n_4529, n_18759);
  or g38926 (n_18861, n_13931, wc196);
  not gc196 (wc196, n_4239);
  nand g38927 (n_14189, n_18750, n_13817);
  nand g38928 (n_18858, n_13931, n_18857);
  nand g38929 (n_20618, n_13931, n_4239);
  or g38930 (n_20619, n_13931, n_4239);
  nand g38931 (n_2033, n_20618, n_20619);
  or g38932 (n_20620, wc197, result[3]);
  not gc197 (wc197, result[5]);
  or g38933 (n_20621, result[5], wc198);
  not gc198 (wc198, result[3]);
  nand g38934 (n_13915, n_20620, n_20621);
  or g38935 (n_19047, wc199, n_19045);
  not gc199 (wc199, n_19044);
  or g38936 (n_18852, wc200, n_3637);
  not gc200 (wc200, n_4528);
  or g38937 (n_18857, n_4240, wc201);
  not gc201 (wc201, n_13439);
  or g38938 (n_18716, n_12774, wc202);
  not gc202 (wc202, result[5]);
  or g38939 (n_18680, n_12765, wc203);
  not gc203 (wc203, result[5]);
  or g38940 (n_18750, n_3637, wc204);
  not gc204 (wc204, n_12553);
  or g38941 (n_18686, n_12766, wc205);
  not gc205 (wc205, result[5]);
  or g38942 (n_18759, n_12764, n_12553);
  or g38943 (n_18692, n_12767, wc206);
  not gc206 (wc206, result[5]);
  nand g38944 (n_18784, n_18779, n_18780);
  or g38945 (n_18722, n_12775, wc207);
  not gc207 (wc207, result[5]);
  or g38946 (n_18698, n_12768, wc208);
  not gc208 (wc208, result[5]);
  nand g38947 (n_18747, n_14463, n_4530);
  or g38948 (n_18704, n_12769, wc209);
  not gc209 (wc209, result[5]);
  nand g38949 (n_18840, n_13439, n_18839);
  or g38950 (n_18710, n_12772, wc210);
  not gc210 (wc210, result[5]);
  nand g38951 (n_4528, n_12860, n_18732);
  nand g38952 (n_20622, n_12860, n_4495);
  or g38953 (n_20623, n_12860, n_4495);
  nand g38954 (n_13782, n_20622, n_20623);
  or g38955 (result[5], n_18674, n_18675);
  nand g38956 (n_18779, n_14497, n_4634);
  nand g38957 (n_12553, n_18737, n_18738);
  nand g38958 (n_18839, n_13945, n_13147);
  or g38959 (n_18746, n_18745, n_12764);
  nand g38960 (n_19045, n_19040, n_19041);
  nand g38961 (n_14463, n_13817, n_18729);
  or g38962 (n_13147, n_11331, n_19602);
  or g38963 (n_18745, wc211, n_4530);
  not gc211 (wc211, n_13828);
  nand g38964 (n_18732, n_13960, n_4496);
  or g38965 (n_19040, wc212, n_13450);
  not gc212 (wc212, n_14469);
  or g38966 (n_18843, n_3637, wc213);
  not gc213 (wc213, n_4529);
  nand g38967 (n_18737, n_14471, n_4530);
  or g38968 (n_18729, n_13828, n_12764);
  or g38969 (n_18675, wc214, n_18673);
  not gc214 (wc214, n_18672);
  or g38970 (n_14497, n_3684, wc215);
  not gc215 (wc215, n_12785);
  or g38971 (n_18758, wc216, n_3637);
  not gc216 (wc216, n_14500);
  nand g38972 (n_4529, n_13960, n_18648);
  or g38973 (n_4496, n_18528, wc217);
  not gc217 (wc217, n_12904);
  nand g38974 (n_5483, n_18569, n_18570);
  nand g38975 (n_5267, n_18593, n_18594);
  or g38976 (n_18738, \data_stack_mem[8] [7], wc218);
  not gc218 (wc218, n_12571);
  nand g38977 (n_5339, n_18563, n_18564);
  nand g38978 (n_20624, \data_stack_mem[8] [7], n_12571);
  or g38979 (n_20625, \data_stack_mem[8] [7], n_12571);
  nand g38980 (n_13828, n_20624, n_20625);
  nand g38981 (n_5051, n_18575, n_18576);
  nand g38982 (n_5411, n_18587, n_18588);
  nand g38983 (n_5555, n_18605, n_18606);
  nand g38984 (n_19602, n_19601, n_18726);
  nand g38985 (n_20626, n_11985, n_11986);
  or g38986 (n_20627, n_11985, n_11986);
  nand g38987 (n_14469, n_20626, n_20627);
  nand g38988 (n_18673, n_18668, n_18669);
  or g38989 (n_18780, wc219, n_12764);
  not gc219 (wc219, n_14496);
  nand g38990 (n_5195, n_18599, n_18600);
  or g38991 (n_20628, result[0], n_13773);
  nand g38992 (n_20629, result[0], n_13773);
  nand g38993 (n_13909, n_20628, n_20629);
  nand g38994 (n_5123, n_18581, n_18582);
  or g38995 (n_12785, n_18642, n_3634);
  or g38996 (n_14500, n_18621, wc220);
  not gc220 (wc220, n_13142);
  nand g38997 (n_12571, n_18615, n_19596);
  nand g38998 (n_18528, n_12905, n_18527);
  or g38999 (n_18599, n_12774, wc221);
  not gc221 (wc221, result[4]);
  or g39000 (n_18569, n_12766, wc222);
  not gc222 (wc222, result[4]);
  or g39004 (n_18593, n_12772, wc223);
  not gc223 (wc223, result[4]);
  nand g39005 (n_4530, n_18626, n_18627);
  nand g39006 (n_11986, n_14277, n_18726);
  or g39007 (n_20632, wc224, result[4]);
  not gc224 (wc224, result[2]);
  or g39008 (n_20633, result[2], wc225);
  not gc225 (wc225, result[4]);
  nand g39009 (n_13773, n_20632, n_20633);
  nand g39010 (n_20634, n_12568, n_12569);
  or g39011 (n_20635, n_12568, n_12569);
  nand g39012 (n_14496, n_20634, n_20635);
  or g39013 (n_18587, n_12769, wc226);
  not gc226 (wc226, result[4]);
  or g39014 (n_18563, n_12765, wc227);
  not gc227 (wc227, result[4]);
  or g39015 (n_18621, n_18620, wc228);
  not gc228 (wc228, n_13146);
  or g39016 (n_18581, n_12768, wc229);
  not gc229 (wc229, result[4]);
  or g39017 (n_18575, n_12767, wc230);
  not gc230 (wc230, result[4]);
  nand g39018 (n_18642, n_18640, n_18641);
  nand g39019 (n_18648, n_4497, n_13146);
  or g39020 (n_19601, wc231, n_11985);
  not gc231 (wc231, n_14277);
  or g39021 (n_18605, n_12775, wc232);
  not gc232 (wc232, result[4]);
  nand g39022 (n_18668, n_14514, n_4634);
  or g39023 (n_20636, wc233, n_4426);
  not gc233 (wc233, n_13908);
  or g39024 (n_20637, n_13908, wc234);
  not gc234 (wc234, n_4426);
  nand g39025 (n_4495, n_20636, n_20637);
  nand g39026 (n_18527, n_14494, n_4432);
  nand g39027 (n_18785, n_18781, n_18782);
  or g39028 (n_19043, n_13996, wc235);
  not gc235 (wc235, n_4242);
  nand g39029 (n_13945, n_13827, n_18645);
  nand g39030 (n_20638, n_13827, n_4208);
  or g39031 (n_20639, n_13827, n_4208);
  nand g39032 (n_4240, n_20638, n_20639);
  or g39033 (n_13146, n_13962, wc236);
  not gc236 (wc236, n_18531);
  or g39034 (n_18640, wc237, n_14070);
  not gc237 (wc237, n_4243);
  or g39035 (n_18641, n_4243, wc238);
  not gc238 (wc238, n_14070);
  or g39036 (n_14514, wc239, n_3693);
  not gc239 (wc239, n_12786);
  nand g39037 (n_5263, n_18467, n_18468);
  nand g39038 (n_12569, n_14272, n_18615);
  nand g39039 (n_5551, n_18479, n_18480);
  nand g39040 (n_5191, n_18473, n_18474);
  or g39041 (n_18627, wc240, n_14483);
  not gc240 (wc240, n_4498);
  nand g39042 (n_5335, n_18437, n_18438);
  or g39043 (result[4], n_18557, n_18558);
  or g39044 (n_18626, n_4498, wc241);
  not gc241 (wc241, n_14483);
  nand g39045 (n_5479, n_18443, n_18444);
  nand g39046 (n_5047, n_18449, n_18450);
  nand g39047 (n_5119, n_18455, n_18456);
  nand g39048 (n_5407, n_18461, n_18462);
  nand g39049 (n_19596, n_14272, n_12568);
  or g39050 (n_18726, \data_stack_mem[8] [7], n_4242);
  or g39051 (n_18479, n_12775, wc242);
  not gc242 (wc242, result[3]);
  nand g39054 (n_13908, n_12904, n_12905);
  or g39055 (n_18473, n_12774, wc243);
  not gc243 (wc243, result[3]);
  or g39056 (n_18461, n_12769, wc244);
  not gc244 (wc244, result[3]);
  or g39057 (n_18645, n_4209, wc245);
  not gc245 (wc245, n_13203);
  or g39058 (n_18467, n_12772, wc246);
  not gc246 (wc246, result[3]);
  nand g39059 (n_18557, n_18553, n_18554);
  nand g39060 (n_18531, n_4498, n_14278);
  nand g39061 (n_11985, n_18611, n_19593);
  nand g39062 (n_4242, n_18632, n_18633);
  or g39063 (n_18455, n_12768, wc247);
  not gc247 (wc247, result[3]);
  nand g39064 (n_14494, n_18402, n_19584);
  nand g39065 (n_14483, n_18500, n_18501);
  or g39066 (n_18449, n_12767, wc248);
  not gc248 (wc248, result[3]);
  nand g39067 (n_13962, data_stack_pointer[3], n_18507);
  or g39068 (n_14070, n_11331, n_18612);
  or g39069 (n_18443, n_12766, wc249);
  not gc249 (wc249, result[3]);
  or g39070 (n_12786, n_18519, n_3634);
  or g39071 (n_18437, n_12765, wc250);
  not gc250 (wc250, result[3]);
  or g39072 (n_18615, \data_stack_mem[8] [6], wc251);
  not gc251 (wc251, n_4531);
  or g39073 (n_18781, wc252, n_14135);
  not gc252 (wc252, n_4531);
  or g39074 (n_18669, wc253, n_12764);
  not gc253 (wc253, n_14513);
  or g39075 (n_13203, n_13957, wc254);
  not gc254 (wc254, n_18522);
  or g39076 (n_12904, n_13142, n_18510);
  nand g39077 (n_18612, n_14264, n_18611);
  nand g39078 (n_18553, n_4634, n_3703);
  or g39079 (n_18500, n_14127, n_12472);
  or g39080 (result[3], n_18431, n_18432);
  nand g39081 (n_12568, n_18489, n_19590);
  or g39082 (n_18501, n_13401, wc255);
  not gc255 (wc255, n_12472);
  nand g39083 (n_20642, n_14058, n_4466);
  or g39084 (n_20643, n_14058, n_4466);
  nand g39085 (n_4498, n_20642, n_20643);
  nand g39086 (n_20644, n_13785, n_13142);
  or g39087 (n_20645, n_13785, n_13142);
  nand g39088 (n_4497, n_20644, n_20645);
  or g39089 (n_18507, \data_stack_mem[7] [7], wc256);
  not gc256 (wc256, n_12472);
  nand g39090 (n_19584, n_13936, n_13142);
  nand g39091 (n_20646, n_14109, n_4499);
  or g39092 (n_20647, n_14109, n_4499);
  nand g39093 (n_4531, n_20646, n_20647);
  nand g39094 (n_18519, n_18517, n_18518);
  nand g39095 (n_20648, n_12566, n_12567);
  or g39096 (n_20649, n_12566, n_12567);
  nand g39097 (n_14513, n_20648, n_20649);
  or g39098 (n_18633, wc257, n_14473);
  not gc257 (wc257, n_4210);
  or g39099 (n_18632, n_4210, wc258);
  not gc258 (wc258, n_14473);
  nand g39100 (n_19593, n_4243, n_14264);
  nand g39104 (n_12472, n_18392, n_19578);
  or g39105 (n_3703, wc259, n_13191);
  not gc259 (wc259, n_14518);
  nand g39106 (n_19590, n_12566, n_14271);
  or g39107 (n_18510, n_13785, n_4432);
  or g39108 (n_14109, n_18393, wc260);
  not gc260 (wc260, data_stack_pointer[3]);
  nand g39109 (n_12567, n_14271, n_18489);
  nand g39110 (n_18611, \data_stack_mem[8] [6], n_11982);
  nand g39111 (n_14473, n_18494, n_18495);
  or g39112 (n_18518, n_4244, wc261);
  not gc261 (wc261, n_14055);
  or g39113 (n_18517, wc262, n_14055);
  not gc262 (wc262, n_4244);
  nand g39114 (n_13957, data_stack_pointer[3], n_18504);
  nand g39115 (n_18674, n_18670, n_18671);
  or g39116 (n_18522, n_4210, wc263);
  not gc263 (wc263, n_14275);
  or g39117 (n_13142, n_14295, wc264);
  not gc264 (wc264, n_18405);
  or g39118 (n_18432, wc265, n_18430);
  not gc265 (wc265, n_18429);
  nand g39119 (n_20652, n_13914, n_4176);
  or g39120 (n_20653, n_13914, n_4176);
  nand g39121 (n_4208, n_20652, n_20653);
  or g39122 (n_18494, n_13401, n_11884);
  or g39123 (n_18495, n_14127, wc266);
  not gc266 (wc266, n_11884);
  nand g39124 (n_18405, n_4466, n_14254);
  nand g39125 (n_20654, n_14060, n_4178);
  or g39126 (n_20655, n_14060, n_4178);
  nand g39127 (n_4210, n_20654, n_20655);
  or g39128 (n_18670, wc267, n_14135);
  not gc267 (wc267, n_4532);
  or g39129 (n_18504, \data_stack_mem[7] [7], n_11884);
  or g39130 (n_14055, n_11331, n_18486);
  nand g39131 (n_13785, n_13936, n_18402);
  nand g39132 (n_11982, n_18485, n_19587);
  nand g39133 (n_20656, n_14016, n_4211);
  or g39134 (n_20657, n_14016, n_4211);
  nand g39135 (n_4243, n_20656, n_20657);
  or g39136 (n_14295, wc268, n_3910);
  not gc268 (wc268, n_18384);
  nand g39137 (n_20658, n_13197, n_4177);
  or g39138 (n_20659, n_13197, n_4177);
  nand g39139 (n_4209, n_20658, n_20659);
  nand g39140 (n_18393, n_14255, n_18392);
  or g39141 (n_18489, \data_stack_mem[8] [5], wc269);
  not gc269 (wc269, n_4532);
  or g39142 (n_18558, wc270, n_18556);
  not gc270 (wc270, n_18555);
  or g39143 (n_13191, wc271, n_3699);
  not gc271 (wc271, n_14517);
  nand g39144 (n_19578, n_4499, n_14255);
  nand g39145 (n_18430, n_18425, n_18426);
  nand g39146 (n_20660, n_14023, n_4467);
  or g39147 (n_20661, n_14023, n_4467);
  nand g39148 (n_4499, n_20660, n_20661);
  nand g39149 (n_18556, n_18551, n_18552);
  nand g39150 (n_20662, n_14114, n_4500);
  or g39151 (n_20663, n_14114, n_4500);
  nand g39152 (n_4532, n_20662, n_20663);
  nand g39153 (n_20664, n_14045, n_4434);
  or g39154 (n_20665, n_14045, n_4434);
  nand g39155 (n_4466, n_20664, n_20665);
  nand g39156 (n_18486, n_14229, n_18485);
  nand g39157 (n_18425, n_14534, n_4634);
  nand g39158 (n_18402, n_13141, n_4433);
  nand g39159 (n_3699, n_18380, n_18381);
  or g39160 (n_18392, \data_stack_mem[7] [6], wc272);
  not gc272 (wc272, n_12469);
  or g39161 (n_18620, n_4426, wc273);
  not gc273 (wc273, n_13141);
  or g39162 (n_18384, \data_stack_mem[6] [7], wc274);
  not gc274 (wc274, n_12373);
  nand g39163 (n_19587, n_4244, n_14229);
  nand g39164 (n_12566, n_18287, n_18288);
  or g39165 (n_13197, n_14228, wc275);
  not gc275 (wc275, n_18387);
  nand g39166 (n_11884, n_18398, n_19581);
  nand g39169 (n_4175, n_14181, n_14257);
  or g39170 (n_14016, n_18399, wc276);
  not gc276 (wc276, data_stack_pointer[3]);
  nand g39171 (n_5547, n_18368, n_18369);
  nand g39172 (n_5043, n_18338, n_18339);
  or g39173 (n_18387, n_4178, wc277);
  not gc277 (wc277, n_14253);
  nand g39174 (n_18287, n_14501, n_12537);
  or g39175 (n_14534, n_3711, wc278);
  not gc278 (wc278, n_12782);
  nand g39176 (n_5115, n_18344, n_18345);
  nand g39177 (n_18399, n_14252, n_18398);
  nand g39178 (n_19581, n_4211, n_14252);
  or g39179 (n_14023, n_18264, n_3910);
  nand g39180 (n_5403, n_18350, n_18351);
  nand g39181 (n_20668, n_13822, n_4144);
  or g39182 (n_20669, n_13822, n_4144);
  nand g39183 (n_4176, n_20668, n_20669);
  or g39184 (n_13141, n_14280, wc279);
  not gc279 (wc279, n_18294);
  nand g39185 (n_12373, n_18263, n_19566);
  or g39186 (n_14114, n_18270, wc280);
  not gc280 (wc280, data_stack_pointer[3]);
  nand g39187 (n_5259, n_18356, n_18357);
  nand g39188 (n_12469, n_18269, n_19569);
  or g39189 (n_14228, wc281, n_3910);
  not gc281 (wc281, n_18282);
  nand g39190 (n_5187, n_18362, n_18363);
  or g39191 (n_18380, n_18379, n_12764);
  nand g39192 (n_5331, n_18326, n_18327);
  or g39193 (n_18551, wc282, n_13450);
  not gc282 (wc282, n_14520);
  nand g39194 (n_18485, \data_stack_mem[8] [5], n_11980);
  nand g39195 (n_5475, n_18332, n_18333);
  or g39196 (n_18288, \data_stack_mem[8] [4], wc283);
  not gc283 (wc283, n_4533);
  nand g39197 (n_20670, n_14024, n_4212);
  or g39198 (n_20671, n_14024, n_4212);
  nand g39199 (n_4244, n_20670, n_20671);
  or g39200 (n_18379, wc284, n_4533);
  not gc284 (wc284, n_13826);
  nand g39201 (n_19569, n_4500, n_14250);
  or g39202 (n_12782, n_18258, n_3634);
  or g39203 (n_18326, n_12765, wc285);
  not gc285 (wc285, result[2]);
  or g39204 (n_18332, n_12766, wc286);
  not gc286 (wc286, result[2]);
  or g39205 (n_18350, n_12769, wc287);
  not gc287 (wc287, result[2]);
  nand g39206 (n_20672, n_13972, n_4400);
  or g39207 (n_20673, n_13972, n_4400);
  nand g39208 (n_4432, n_20672, n_20673);
  or g39209 (n_18338, n_12767, wc288);
  not gc288 (wc288, result[2]);
  or g39210 (n_18282, \data_stack_mem[6] [7], n_11783);
  nand g39211 (n_4433, n_13972, n_18291);
  or g39212 (n_18356, n_12772, wc289);
  not gc289 (wc289, result[2]);
  or g39213 (n_18362, n_12774, wc290);
  not gc290 (wc290, result[2]);
  nand g39214 (n_20674, n_13220, n_4145);
  or g39215 (n_20675, n_13220, n_4145);
  nand g39216 (n_4177, n_20674, n_20675);
  nand g39217 (n_18270, n_14250, n_18269);
  or g39218 (n_18368, n_12775, wc291);
  not gc291 (wc291, result[2]);
  or g39219 (n_14280, n_3908, wc292);
  not gc292 (wc292, n_18237);
  nand g39220 (n_20676, n_14030, n_4146);
  or g39221 (n_20677, n_14030, n_4146);
  nand g39222 (n_4178, n_20676, n_20677);
  or g39223 (n_18344, n_12768, wc293);
  not gc293 (wc293, result[2]);
  nand g39224 (n_18264, n_14304, n_18263);
  nand g39225 (n_18381, n_14515, n_4533);
  nand g39226 (n_18294, n_4434, n_14305);
  nand g39227 (n_18398, \data_stack_mem[7] [6], n_11881);
  nand g39228 (n_19566, n_4467, n_14304);
  nand g39229 (n_11980, n_18372, n_19575);
  nand g39230 (n_20678, n_11944, n_11978);
  or g39231 (n_20679, n_11944, n_11978);
  nand g39232 (n_14520, n_20678, n_20679);
  or g39233 (n_4426, n_18243, wc294);
  not gc294 (wc294, n_12814);
  nand g39234 (n_11881, n_18275, n_19572);
  or g39235 (n_13220, n_14300, wc295);
  not gc295 (wc295, n_18240);
  nand g39236 (n_20680, n_14000, n_4179);
  or g39237 (n_20681, n_14000, n_4179);
  nand g39238 (n_4211, n_20680, n_20681);
  or g39239 (n_18237, \data_stack_mem[5] [7], wc296);
  not gc296 (wc296, n_12274);
  nand g39240 (n_18258, n_18256, n_18257);
  nand g39241 (n_11783, n_18233, n_19563);
  or g39242 (n_18269, \data_stack_mem[7] [5], wc297);
  not gc297 (wc297, n_12467);
  nand g39243 (n_11978, n_14262, n_18372);
  nand g39244 (n_20682, n_14039, n_4435);
  or g39245 (n_20683, n_14039, n_4435);
  nand g39246 (n_4467, n_20682, n_20683);
  nand g39247 (n_20684, n_14038, n_4402);
  or g39248 (n_20685, n_14038, n_4402);
  nand g39249 (n_4434, n_20684, n_20685);
  nand g39250 (n_19575, n_14262, n_11944);
  or g39251 (n_4533, wc298, n_18222);
  not gc298 (wc298, n_18221);
  or g39252 (n_14024, n_18276, wc299);
  not gc299 (wc299, data_stack_pointer[3]);
  nand g39253 (n_20686, n_14040, n_4468);
  or g39254 (n_20687, n_14040, n_4468);
  nand g39255 (n_4500, n_20686, n_20687);
  or g39256 (n_18263, \data_stack_mem[6] [6], wc300);
  not gc300 (wc300, n_12370);
  nand g39257 (n_14515, n_13817, n_18279);
  or g39258 (result[2], n_18320, n_18321);
  nand g39259 (n_18291, n_4401, n_12814);
  or g39260 (n_18240, n_4146, wc301);
  not gc301 (wc301, n_14279);
  or g39261 (n_12814, n_14317, wc302);
  not gc302 (wc302, n_18201);
  or g39262 (n_14040, n_18066, n_3910);
  or g39263 (n_14039, n_18183, n_3908);
  or g39264 (n_18257, n_4246, wc303);
  not gc303 (wc303, n_14031);
  nand g39265 (n_12274, n_18182, n_19551);
  nand g39266 (n_5399, n_18158, n_18159);
  nand g39267 (n_19563, n_4179, n_14309);
  nand g39268 (n_5543, n_18176, n_18177);
  nand g39269 (n_18320, n_18316, n_18317);
  nand g39270 (n_5255, n_18164, n_18165);
  or g39271 (n_18279, n_13826, n_12764);
  nand g39272 (n_12370, n_18065, n_19542);
  or g39273 (n_18554, n_13996, wc304);
  not gc304 (wc304, n_4245);
  nand g39274 (n_5327, n_18134, n_18135);
  nand g39275 (n_5183, n_18170, n_18171);
  nand g39276 (n_5111, n_18152, n_18153);
  nand g39277 (n_18276, n_14261, n_18275);
  nand g39278 (n_19572, n_4212, n_14261);
  or g39279 (n_18256, wc305, n_14031);
  not gc305 (wc305, n_4246);
  or g39280 (n_14000, n_18234, n_3910);
  nand g39281 (n_18222, n_18219, n_18220);
  nand g39282 (n_18372, \data_stack_mem[8] [4], n_4245);
  nand g39283 (n_5471, n_18140, n_18141);
  nand g39284 (n_12467, n_18206, n_18207);
  nand g39285 (n_5039, n_18146, n_18147);
  nand g39286 (n_20688, n_13809, n_4112);
  or g39287 (n_20689, n_13809, n_4112);
  nand g39288 (n_4144, n_20688, n_20689);
  or g39289 (n_14300, n_3908, wc306);
  not gc306 (wc306, n_18198);
  nand g39290 (n_18201, n_14274, n_4402);
  nand g39291 (n_18183, n_14313, n_18182);
  or g39292 (n_18426, wc307, n_12764);
  not gc307 (wc307, n_14533);
  or g39293 (n_14317, n_20, wc308);
  not gc308 (wc308, n_18096);
  nand g39294 (n_18317, n_4634, n_3721);
  or g39295 (n_18134, n_12765, wc309);
  not gc309 (wc309, result[1]);
  nand g39296 (n_19551, n_4435, n_14313);
  nand g39297 (n_18275, \data_stack_mem[7] [5], n_11879);
  or g39298 (n_18198, \data_stack_mem[5] [7], n_11682);
  nand g39299 (n_18234, n_14309, n_18233);
  or g39300 (n_18140, n_12766, wc310);
  not gc310 (wc310, result[1]);
  nand g39301 (n_20690, n_12813, n_4113);
  or g39302 (n_20691, n_12813, n_4113);
  nand g39303 (n_4145, n_20690, n_20691);
  or g39304 (n_18146, n_12767, wc311);
  not gc311 (wc311, result[1]);
  nand g39305 (n_20692, n_14035, n_4147);
  or g39306 (n_20693, n_14035, n_4147);
  nand g39307 (n_4179, n_20692, n_20693);
  nand g39308 (n_18066, n_14314, n_18065);
  or g39309 (n_18158, n_12769, wc312);
  not gc312 (wc312, result[1]);
  or g39310 (n_18321, wc313, n_18319);
  not gc313 (wc313, n_18318);
  or g39311 (n_18164, n_12772, wc314);
  not gc314 (wc314, result[1]);
  or g39312 (n_18170, n_12774, wc315);
  not gc315 (wc315, result[1]);
  nand g39313 (n_20694, \data_stack_mem[8] [4], n_12537);
  or g39314 (n_20695, \data_stack_mem[8] [4], n_12537);
  nand g39315 (n_13826, n_20694, n_20695);
  nand g39316 (n_19542, n_4468, n_14314);
  or g39317 (n_14031, n_11331, n_18228);
  nand g39318 (n_4245, n_18248, n_18249);
  or g39319 (n_18176, n_12775, wc316);
  not gc316 (wc316, result[1]);
  or g39320 (n_18219, n_14145, n_14283);
  or g39321 (n_18206, \data_stack_mem[7] [4], wc317);
  not gc317 (wc317, n_14283);
  or g39322 (n_18220, n_18218, wc318);
  not gc318 (wc318, n_12438);
  nand g39323 (n_11944, n_18227, n_19560);
  nand g39324 (n_20696, n_14085, n_4114);
  or g39325 (n_20697, n_14085, n_4114);
  nand g39326 (n_4146, n_20696, n_20697);
  or g39327 (n_18152, n_12768, wc319);
  not gc319 (wc319, result[1]);
  or g39328 (n_18065, \data_stack_mem[6] [5], wc320);
  not gc320 (wc320, n_12368);
  or g39329 (n_12813, n_14286, wc321);
  not gc321 (wc321, n_18093);
  nand g39330 (n_12537, n_18186, n_19554);
  nand g39331 (n_19560, n_4246, n_14287);
  nand g39332 (n_18233, \data_stack_mem[6] [6], n_11780);
  or g39333 (n_18218, n_4501, n_13403);
  nand g39334 (n_18207, n_4501, n_12438);
  nand g39335 (n_18221, n_14502, n_4501);
  nand g39336 (n_20698, n_14036, n_4436);
  or g39337 (n_20699, n_14036, n_4436);
  nand g39338 (n_4468, n_20698, n_20699);
  nand g39339 (n_4401, n_13906, n_18195);
  or g39340 (n_18249, wc322, n_14489);
  not gc322 (wc322, n_4213);
  nand g39341 (n_18228, n_14287, n_18227);
  or g39342 (n_18248, n_4213, wc323);
  not gc323 (wc323, n_14489);
  nand g39343 (n_18319, n_18314, n_18315);
  nand g39344 (n_20700, n_14032, n_4403);
  or g39345 (n_20701, n_14032, n_4403);
  nand g39346 (n_4435, n_20700, n_20701);
  nand g39347 (n_20702, n_14043, n_4180);
  or g39348 (n_20703, n_14043, n_4180);
  nand g39349 (n_4212, n_20702, n_20703);
  nand g39350 (n_11682, n_18071, n_19545);
  nand g39351 (n_11879, n_18191, n_19557);
  or g39352 (n_18096, \data_stack_mem[4] [7], wc324);
  not gc324 (wc324, n_12175);
  or g39353 (n_3721, wc325, n_13189);
  not gc325 (wc325, n_14538);
  nand g39354 (n_20704, n_13941, n_13906);
  or g39355 (n_20705, n_13941, n_13906);
  nand g39356 (n_4400, n_20704, n_20705);
  or g39357 (result[1], n_18128, n_18129);
  nand g39358 (n_20706, n_12562, n_12563);
  or g39359 (n_20707, n_12562, n_12563);
  nand g39360 (n_14533, n_20706, n_20707);
  or g39361 (n_14035, n_18072, n_3908);
  or g39362 (n_18182, \data_stack_mem[5] [6], wc326);
  not gc326 (wc326, n_12271);
  nand g39363 (n_4402, n_18101, n_18102);
  nand g39364 (n_12175, n_18023, n_19530);
  nand g39365 (n_19545, n_4147, n_14299);
  or g39366 (n_14286, n_20, wc327);
  not gc327 (wc327, n_18048);
  nand g39367 (n_18431, n_18427, n_18428);
  or g39368 (n_18243, wc328, n_13941);
  not gc328 (wc328, n_12809);
  or g39369 (n_14036, n_18030, n_3908);
  or g39370 (n_14502, n_18045, wc329);
  not gc329 (wc329, data_stack_pointer[3]);
  nand g39371 (n_19554, n_12562, n_14259);
  nand g39372 (n_18128, n_18124, n_18125);
  or g39373 (n_18093, wc330, n_4114);
  not gc330 (wc330, n_14316);
  nand g39374 (n_12368, n_17969, n_19515);
  nand g39375 (n_11780, n_18077, n_19548);
  nand g39376 (n_18227, \data_stack_mem[8] [3], n_11976);
  nand g39377 (n_12271, n_18029, n_19533);
  nand g39378 (n_18195, n_4369, n_12809);
  nand g39381 (n_4112, n_13928, n_14063);
  or g39382 (n_14032, n_20, n_18024);
  nand g39383 (n_14489, n_18083, n_18084);
  or g39384 (n_18314, wc331, n_13450);
  not gc331 (wc331, n_14540);
  or g39385 (n_14043, n_18078, n_3910);
  nand g39386 (n_19557, n_4213, n_14307);
  or g39387 (n_13189, wc332, n_3717);
  not gc332 (wc332, n_14537);
  nand g39388 (n_12563, n_14259, n_18186);
  nand g39389 (n_18072, n_14299, n_18071);
  nand g39390 (n_20710, n_14014, n_4469);
  or g39391 (n_20711, n_14014, n_4469);
  nand g39392 (n_4501, n_20710, n_20711);
  or g39393 (n_18048, \data_stack_mem[4] [7], n_11581);
  nand g39394 (n_19515, n_4469, n_14268);
  nand g39395 (n_5395, n_17945, n_17946);
  nand g39396 (n_18071, \data_stack_mem[5] [6], n_11679);
  or g39397 (n_18427, wc333, n_14135);
  not gc333 (wc333, n_4534);
  nand g39398 (n_19548, n_4180, n_14310);
  nand g39399 (n_18030, n_14256, n_18029);
  nand g39400 (n_3717, n_18089, n_18090);
  nand g39401 (n_20712, n_14013, n_4214);
  or g39402 (n_20713, n_14013, n_4214);
  nand g39403 (n_4246, n_20712, n_20713);
  nand g39404 (n_5323, n_17921, n_17922);
  or g39405 (n_14014, n_17970, n_3910);
  nand g39406 (n_11976, n_18060, n_19539);
  nand g39407 (n_5179, n_17951, n_17952);
  nand g39408 (n_5467, n_17927, n_17928);
  nand g39409 (n_4114, n_18053, n_18054);
  or g39410 (n_18084, n_14145, wc334);
  not gc334 (wc334, n_11843);
  or g39411 (n_12809, n_13943, wc335);
  not gc335 (wc335, n_18057);
  or g39412 (n_18083, n_13403, n_11843);
  nand g39413 (n_18078, n_14310, n_18077);
  or g39414 (n_18102, wc336, n_14510);
  not gc336 (wc336, n_4370);
  nand g39415 (n_18045, n_18043, n_18044);
  nand g39416 (n_5251, n_17957, n_17958);
  nand g39417 (n_19530, n_4403, n_14247);
  nand g39418 (n_5035, n_17933, n_17934);
  nand g39419 (n_20714, n_14011, n_4115);
  or g39420 (n_20715, n_14011, n_4115);
  nand g39421 (n_4147, n_20714, n_20715);
  nand g39422 (n_18191, \data_stack_mem[7] [4], n_11843);
  or g39423 (n_18101, n_4370, wc337);
  not gc337 (wc337, n_14510);
  nand g39424 (n_5107, n_17939, n_17940);
  nand g39425 (n_20716, n_11925, n_11974);
  or g39426 (n_20717, n_11925, n_11974);
  nand g39427 (n_14540, n_20716, n_20717);
  nand g39428 (n_5539, n_17963, n_17964);
  nand g39429 (n_20718, n_12824, n_4081);
  or g39430 (n_20719, n_12824, n_4081);
  nand g39431 (n_4113, n_20718, n_20719);
  or g39432 (n_18129, wc338, n_18127);
  not gc338 (wc338, n_18126);
  or g39433 (n_18186, \data_stack_mem[8] [3], wc339);
  not gc339 (wc339, n_4534);
  nand g39434 (n_18024, n_14247, n_18023);
  nand g39435 (n_19533, n_4436, n_14256);
  nand g39436 (n_18125, n_4634, n_3730);
  or g39437 (n_18023, \data_stack_mem[4] [6], wc340);
  not gc340 (wc340, n_12172);
  or g39438 (n_17927, n_12766, result[0]);
  nand g39439 (n_20720, n_14025, n_4502);
  or g39440 (n_20721, n_14025, n_4502);
  nand g39441 (n_4534, n_20720, n_20721);
  nand g39442 (n_18077, \data_stack_mem[6] [5], n_11778);
  or g39443 (n_17921, n_12765, result[0]);
  nand g39444 (n_14510, n_17999, n_18000);
  or g39445 (n_17933, n_12767, result[0]);
  or g39446 (n_14011, n_20, n_17988);
  or g39447 (n_18044, wc341, n_12438);
  not gc341 (wc341, \data_stack_mem[7] [4]);
  or g39448 (n_17939, n_12768, result[0]);
  nand g39449 (n_11679, n_17981, n_19521);
  or g39450 (n_18043, \data_stack_mem[7] [4], wc342);
  not gc342 (wc342, n_12438);
  nand g39451 (n_18057, n_4370, n_14315);
  nand g39452 (n_20722, n_14009, n_4148);
  or g39453 (n_20723, n_14009, n_4148);
  nand g39454 (n_4180, n_20722, n_20723);
  or g39455 (n_17945, n_12769, result[0]);
  nand g39456 (n_17970, n_14268, n_17969);
  or g39457 (n_17951, n_12774, result[0]);
  nand g39458 (n_20724, n_14089, n_4437);
  or g39459 (n_20725, n_14089, n_4437);
  nand g39460 (n_4469, n_20724, n_20725);
  nand g39461 (n_11843, n_18035, n_19536);
  or g39462 (n_18089, wc343, n_12764);
  not gc343 (wc343, n_14535);
  nand g39463 (n_13943, n_37, n_18003);
  nand g39464 (n_18127, n_18122, n_18123);
  nand g39465 (n_11581, n_17987, n_19524);
  nand g39466 (n_20726, n_14012, n_4181);
  or g39467 (n_20727, n_14012, n_4181);
  nand g39468 (n_4213, n_20726, n_20727);
  or g39469 (n_3730, wc344, n_13233);
  not gc344 (wc344, n_14552);
  or g39470 (n_18029, \data_stack_mem[5] [5], wc345);
  not gc345 (wc345, n_12269);
  or g39471 (n_18053, n_4082, wc346);
  not gc346 (wc346, n_14506);
  or g39472 (n_18054, wc347, n_14506);
  not gc347 (wc347, n_4082);
  or g39473 (n_14013, n_18036, wc348);
  not gc348 (wc348, data_stack_pointer[3]);
  nand g39474 (n_20728, n_14098, n_4404);
  or g39475 (n_20729, n_14098, n_4404);
  nand g39476 (n_4436, n_20728, n_20729);
  nand g39477 (n_19539, n_14298, n_11925);
  or g39478 (n_12824, n_13944, wc349);
  not gc349 (wc349, n_18006);
  nand g39479 (n_11974, n_14298, n_18060);
  or g39480 (n_17963, n_12775, result[0]);
  or g39481 (n_17957, n_12772, result[0]);
  nand g39482 (n_12438, n_17975, n_19518);
  or g39483 (n_18122, wc350, n_13450);
  not gc350 (wc350, n_14554);
  or g39484 (n_18006, n_4082, wc351);
  not gc351 (wc351, n_14248);
  nand g39485 (n_18036, n_14282, n_18035);
  or g39486 (n_14098, n_20, n_17877);
  nand g39487 (n_13944, n_37, n_17910);
  nand g39488 (n_12269, n_17801, n_19482);
  nand g39489 (n_18060, \data_stack_mem[8] [2], n_4247);
  nand g39490 (n_14506, n_17897, n_17898);
  or g39491 (n_18003, \data_stack_mem[3] [7], wc352);
  not gc352 (wc352, n_12079);
  or g39492 (n_20730, wc353, n_13818);
  not gc353 (wc353, n_12515);
  or g39493 (n_20731, n_12515, wc354);
  not gc354 (wc354, n_13818);
  nand g39494 (n_14535, n_20730, n_20731);
  or g39495 (n_14012, n_17994, n_3910);
  or g39496 (n_18316, n_13996, wc355);
  not gc355 (wc355, n_4247);
  nand g39497 (result[0], n_14576, n_4634);
  nand g39498 (n_19524, n_4115, n_14238);
  nand g39499 (n_19521, n_4148, n_14311);
  or g39500 (n_14089, n_17802, n_3908);
  nand g39501 (n_12562, n_18011, n_18012);
  or g39502 (n_17969, \data_stack_mem[6] [4], wc356);
  not gc356 (wc356, n_12339);
  or g39503 (n_14009, n_17982, n_3908);
  nand g39504 (n_19536, n_4214, n_14282);
  or g39505 (n_18000, n_13765, wc357);
  not gc357 (wc357, n_12079);
  or g39506 (n_17999, n_14136, n_12079);
  nand g39507 (n_17988, n_14238, n_17987);
  nand g39508 (n_20732, n_14111, n_4371);
  or g39509 (n_20733, n_14111, n_4371);
  nand g39510 (n_4403, n_20732, n_20733);
  nand g39511 (n_11778, n_17993, n_19527);
  or g39512 (n_13233, wc358, n_3726);
  not gc358 (wc358, n_14551);
  nand g39513 (n_12172, n_17876, n_19503);
  or g39514 (n_14025, n_17976, wc359);
  not gc359 (wc359, data_stack_pointer[3]);
  nand g39515 (n_19503, n_4404, n_14198);
  nand g39516 (n_18035, \data_stack_mem[7] [3], n_11875);
  or g39517 (n_14111, wc360, n_17883);
  not gc360 (wc360, n_37);
  or g39518 (n_20734, wc361, n_11973);
  not gc361 (wc361, n_13921);
  or g39519 (n_20735, n_13921, wc362);
  not gc362 (wc362, n_11973);
  nand g39520 (n_14554, n_20734, n_20735);
  nand g39521 (n_17994, n_14312, n_17993);
  or g39522 (n_14576, wc363, n_17859);
  not gc363 (wc363, n_17858);
  nand g39523 (n_20736, \data_stack_mem[8] [2], n_4535);
  or g39524 (n_20737, \data_stack_mem[8] [2], n_4535);
  nand g39525 (n_13818, n_20736, n_20737);
  nand g39526 (n_4247, n_18017, n_18018);
  or g39527 (n_18090, n_13817, wc364);
  not gc364 (wc364, n_4535);
  nand g39528 (n_19482, n_4437, n_14230);
  nand g39529 (n_11925, n_17886, n_19509);
  nand g39530 (n_17877, n_14198, n_17876);
  nand g39531 (n_19518, n_4502, n_14308);
  nand g39532 (n_12079, n_17882, n_19506);
  or g39533 (n_17910, \data_stack_mem[3] [7], n_11483);
  or g39534 (n_17898, n_14136, wc365);
  not gc365 (wc365, n_11483);
  or g39535 (n_17897, n_13765, n_11483);
  nand g39536 (n_20738, n_14099, n_4116);
  or g39537 (n_20739, n_14099, n_4116);
  nand g39538 (n_4148, n_20738, n_20739);
  nand g39539 (n_17802, n_14230, n_17801);
  nand g39540 (n_12339, n_17807, n_19485);
  nand g39541 (n_20740, n_14102, n_4083);
  or g39542 (n_20741, n_14102, n_4083);
  nand g39543 (n_4115, n_20740, n_20741);
  nand g39544 (n_17982, n_14311, n_17981);
  nand g39545 (n_18011, n_14521, n_4535);
  nand g39546 (n_3726, n_17906, n_17907);
  nand g39547 (n_19527, n_4181, n_14312);
  nand g39548 (n_17987, \data_stack_mem[4] [6], n_11578);
  nand g39549 (n_17976, n_14308, n_17975);
  nand g39550 (n_17883, n_14203, n_17882);
  or g39551 (n_18018, wc366, n_14493);
  not gc366 (wc366, n_4215);
  or g39552 (n_18017, n_4215, wc367);
  not gc367 (wc367, n_14493);
  nand g39553 (n_11578, n_17819, n_19491);
  nand g39554 (n_11483, n_17825, n_19494);
  or g39555 (n_20742, wc368, n_4330);
  not gc368 (wc368, n_12897);
  or g39556 (n_20743, n_12897, wc369);
  not gc369 (wc369, n_4330);
  nand g39557 (n_4369, n_20742, n_20743);
  nand g39558 (n_17859, n_17856, n_17857);
  or g39559 (n_17975, \data_stack_mem[7] [3], wc370);
  not gc370 (wc370, n_12463);
  nand g39560 (n_17981, \data_stack_mem[5] [5], n_11677);
  nand g39561 (n_20744, n_14075, n_4050);
  or g39562 (n_20745, n_14075, n_4050);
  nand g39563 (n_4082, n_20744, n_20745);
  or g39564 (n_17876, \data_stack_mem[4] [5], wc371);
  not gc371 (wc371, n_12170);
  or g39565 (n_17801, \data_stack_mem[5] [4], wc372);
  not gc372 (wc372, n_12240);
  nand g39566 (n_20746, n_13998, n_4182);
  or g39567 (n_20747, n_13998, n_4182);
  nand g39568 (n_4214, n_20746, n_20747);
  or g39569 (n_14102, wc373, n_17826);
  not gc373 (wc373, n_37);
  or g39570 (n_19509, n_13921, wc374);
  not gc374 (wc374, n_14303);
  nand g39571 (n_20748, n_14108, n_4405);
  or g39572 (n_20749, n_14108, n_4405);
  nand g39573 (n_4437, n_20748, n_20749);
  nand g39574 (n_4535, n_17915, n_17916);
  nand g39575 (n_11875, n_17891, n_19512);
  or g39576 (n_18012, \data_stack_mem[8] [2], wc375);
  not gc375 (wc375, n_12515);
  nand g39577 (n_20750, n_14116, n_4338);
  or g39578 (n_20751, n_14116, n_4338);
  nand g39579 (n_4370, n_20750, n_20751);
  nand g39580 (n_19485, n_4470, n_14293);
  nand g39581 (n_13941, n_4330, n_12897);
  nand g39582 (n_19506, n_4371, n_14203);
  or g39583 (n_14099, n_20, n_17820);
  nand g39584 (n_20752, n_14120, n_4470);
  or g39585 (n_20753, n_14120, n_4470);
  nand g39586 (n_4502, n_20752, n_20753);
  nand g39587 (n_20754, n_12895, n_4049);
  or g39588 (n_20755, n_12895, n_4049);
  nand g39589 (n_4081, n_20754, n_20755);
  nand g39590 (n_17907, n_14549, n_4536);
  nand g39591 (n_17993, \data_stack_mem[6] [4], n_11742);
  nand g39592 (n_20756, n_14003, n_4149);
  or g39593 (n_20757, n_14003, n_4149);
  nand g39594 (n_4181, n_20756, n_20757);
  nand g39595 (n_11973, n_14303, n_17886);
  nand g39596 (n_11677, n_17813, n_19488);
  nand g39597 (n_17826, n_14204, n_17825);
  nand g39598 (n_20758, n_14107, n_4438);
  or g39599 (n_20759, n_14107, n_4438);
  nand g39600 (n_4470, n_20758, n_20759);
  or g39601 (n_14003, n_17814, n_3908);
  nand g39602 (n_19494, n_4083, n_14204);
  nand g39603 (n_12463, n_17843, n_19500);
  or g39604 (n_14120, n_17808, n_3910);
  or g39605 (n_12895, n_14219, wc376);
  not gc376 (wc376, n_17865);
  nand g39606 (n_17820, n_14197, n_17819);
  or g39607 (n_14108, n_20, n_17745);
  nand g39608 (n_12240, n_17690, n_19452);
  nand g39609 (n_17857, n_14574, n_625);
  nand g39610 (n_19491, n_4116, n_14197);
  nand g39611 (n_12515, n_17870, n_17871);
  or g39612 (n_17906, n_17905, n_12764);
  nand g39613 (n_19512, n_4215, n_14276);
  or g39614 (n_13998, n_17832, n_3910);
  or g39615 (n_17915, n_4503, wc377);
  not gc377 (wc377, n_14523);
  or g39616 (n_17916, wc378, n_14523);
  not gc378 (wc378, n_4503);
  nand g39617 (n_12170, n_17744, n_19476);
  or g39618 (n_12897, n_14218, wc379);
  not gc379 (wc379, n_17862);
  nand g39619 (n_14493, n_17837, n_17838);
  nand g39620 (n_11742, n_17831, n_19497);
  or g39621 (n_18124, n_13996, wc380);
  not gc380 (wc380, n_4248);
  nand g39622 (n_14549, n_13817, n_17847);
  or g39623 (n_17882, \data_stack_mem[3] [6], wc381);
  not gc381 (wc381, n_12076);
  nand g39624 (n_17886, \data_stack_mem[8] [1], n_4248);
  nand g39625 (n_20760, n_14090, n_4372);
  or g39626 (n_20761, n_14090, n_4372);
  nand g39627 (n_4404, n_20760, n_20761);
  nand g39628 (n_14218, n_3902, n_17766);
  nand g39629 (n_19500, n_4503, n_14260);
  nand g39630 (n_17862, n_14210, n_4338);
  nand g39631 (n_17832, n_14290, n_17831);
  or g39632 (n_14090, wc382, n_17751);
  not gc382 (wc382, n_37);
  nand g39633 (n_14523, n_17762, n_17763);
  or g39634 (n_17847, n_13830, n_12764);
  or g39635 (n_14107, n_17691, n_3908);
  or g39636 (n_17905, wc383, n_4536);
  not gc383 (wc383, n_13830);
  nand g39637 (n_17819, \data_stack_mem[4] [5], n_11576);
  or g39638 (n_4248, wc384, n_17796);
  not gc384 (wc384, n_17795);
  nand g39639 (n_17891, \data_stack_mem[7] [2], n_11824);
  nand g39640 (n_625, n_17756, n_17757);
  nand g39641 (n_19488, n_4149, n_14195);
  nand g39642 (n_19497, n_4182, n_14290);
  nand g39643 (n_19452, n_4438, n_14201);
  nand g39644 (n_17870, n_14527, n_4536);
  nand g39645 (n_17745, n_14207, n_17744);
  nand g39646 (n_12076, n_17750, n_19479);
  nand g39647 (n_17825, \data_stack_mem[3] [6], n_11480);
  nand g39648 (n_14219, n_3902, n_17769);
  nand g39649 (n_20762, n_14113, n_4084);
  or g39650 (n_20763, n_14113, n_4084);
  nand g39651 (n_4116, n_20762, n_20763);
  or g39652 (n_17865, wc385, n_4050);
  not gc385 (wc385, n_14211);
  or g39653 (n_17838, n_14152, wc386);
  not gc386 (wc386, n_11824);
  or g39654 (n_17837, n_13402, n_11824);
  nand g39655 (n_17814, n_14195, n_17813);
  nand g39656 (n_17808, n_14293, n_17807);
  nand g39657 (n_19476, n_14207, n_4405);
  or g39658 (n_17769, \data_stack_mem[2] [7], n_12648);
  nand g39659 (n_11576, n_17708, n_19461);
  nand g39660 (n_20764, n_14110, n_4117);
  or g39661 (n_20765, n_14110, n_4117);
  nand g39662 (n_4149, n_20764, n_20765);
  nand g39663 (n_20766, n_14100, n_4406);
  or g39664 (n_20767, n_14100, n_4406);
  nand g39665 (n_4438, n_20766, n_20767);
  or g39666 (n_17744, \data_stack_mem[4] [4], wc387);
  not gc387 (wc387, n_12141);
  nand g39667 (n_20768, n_14103, n_4051);
  or g39668 (n_20769, n_14103, n_4051);
  nand g39669 (n_4083, n_20768, n_20769);
  nand g39670 (n_17831, \data_stack_mem[6] [3], n_11774);
  nand g39671 (n_19479, n_14214, n_4372);
  nand g39672 (n_17796, n_17793, n_17794);
  nand g39673 (n_11480, n_17714, n_19464);
  or g39674 (n_17757, n_13409, n_11331);
  nand g39675 (n_17691, n_14201, n_17690);
  nand g39676 (n_17795, n_14505, n_4216);
  or g39677 (n_17871, \data_stack_mem[8] [1], wc388);
  not gc388 (wc388, n_13409);
  nand g39678 (n_20770, \data_stack_mem[8] [1], n_13409);
  or g39679 (n_20771, \data_stack_mem[8] [1], n_13409);
  nand g39680 (n_13830, n_20770, n_20771);
  nand g39681 (n_4536, n_17774, n_17775);
  nand g39682 (n_17813, \data_stack_mem[5] [4], n_11641);
  nand g39683 (n_20772, n_14078, n_4339);
  or g39684 (n_20773, n_14078, n_4339);
  nand g39685 (n_4371, n_20772, n_20773);
  nand g39686 (n_17751, n_14214, n_17750);
  nand g39687 (n_20774, n_14084, n_4183);
  or g39688 (n_20775, n_14084, n_4183);
  nand g39689 (n_4215, n_20774, n_20775);
  nand g39690 (n_20776, n_14087, n_4471);
  or g39691 (n_20777, n_14087, n_4471);
  nand g39692 (n_4503, n_20776, n_20777);
  or g39693 (n_17763, n_13402, wc389);
  not gc389 (wc389, n_12416);
  or g39694 (n_17807, \data_stack_mem[6] [3], wc390);
  not gc390 (wc390, n_12364);
  nand g39695 (n_11824, n_17780, n_17781);
  or g39696 (n_14113, wc391, n_17715);
  not gc391 (wc391, n_37);
  or g39697 (n_17843, \data_stack_mem[7] [2], wc392);
  not gc392 (wc392, n_12416);
  or g39698 (n_17762, n_14152, n_12416);
  nand g39699 (n_20778, n_14112, n_4150);
  or g39700 (n_20779, n_14112, n_4150);
  nand g39701 (n_4182, n_20778, n_20779);
  or g39702 (n_17766, \data_stack_mem[2] [7], wc393);
  not gc393 (wc393, n_12725);
  nand g39703 (n_17715, n_14213, n_17714);
  nand g39704 (n_12725, n_17684, n_19449);
  or g39705 (n_17775, wc394, n_14529);
  not gc394 (wc394, n_4504);
  nand g39706 (n_12141, n_17579, n_19419);
  or g39707 (n_17774, n_4504, wc395);
  not gc395 (wc395, n_14529);
  or g39708 (n_17794, n_13400, n_14291);
  or g39709 (n_17793, n_13813, n_17792);
  nand g39710 (n_19464, n_14213, n_4084);
  or g39711 (n_14505, n_17649, wc396);
  not gc396 (wc396, data_stack_pointer[3]);
  or g39712 (n_14087, n_17697, n_3910);
  or g39713 (n_14110, n_20, n_17709);
  nand g39714 (n_12648, n_17720, n_19467);
  or g39715 (n_14078, n_17685, wc397);
  not gc397 (wc397, n_3902);
  or g39716 (n_14103, n_17721, wc398);
  not gc398 (wc398, n_3902);
  nand g39717 (n_4405, n_17738, n_17739);
  or g39718 (n_14084, n_17727, n_3910);
  nand g39719 (n_12416, n_17732, n_19473);
  nand g39720 (n_12364, n_17696, n_19455);
  nand g39721 (n_19461, n_14205, n_4117);
  or g39722 (n_17690, \data_stack_mem[5] [3], wc399);
  not gc399 (wc399, n_12265);
  or g39723 (n_14112, n_17703, n_3908);
  nand g39724 (n_11641, n_17702, n_19458);
  nand g39725 (n_17780, \data_stack_mem[7] [1], n_14291);
  or g39726 (n_14100, n_20, n_17580);
  or g39727 (n_17750, \data_stack_mem[3] [5], wc400);
  not gc400 (wc400, n_12074);
  nand g39728 (n_11774, n_17726, n_19470);
  nand g39729 (n_17756, n_1425, n_14302);
  nand g39730 (n_12074, n_17639, n_19446);
  nand g39731 (n_19419, n_4406, n_14217);
  nand g39732 (n_1425, n_17678, n_17679);
  or g39733 (n_17792, n_4216, n_14151);
  nand g39734 (n_17649, n_17647, n_17648);
  nand g39735 (n_17685, n_14225, n_17684);
  or g39736 (n_17738, n_4373, wc401);
  not gc401 (wc401, n_14491);
  or g39737 (n_17739, wc402, n_14491);
  not gc402 (wc402, n_4373);
  nand g39738 (n_17727, n_14233, n_17726);
  nand g39739 (n_12265, n_17585, n_19422);
  or g39740 (n_17781, n_13813, wc403);
  not gc403 (wc403, n_4216);
  nand g39741 (n_17580, n_14217, n_17579);
  nand g39742 (n_17703, n_14202, n_17702);
  nand g39743 (n_19449, n_4339, n_14225);
  nand g39744 (n_14529, n_17654, n_17655);
  nand g39745 (n_17697, n_14236, n_17696);
  nand g39746 (n_19467, n_4051, n_14224);
  nand g39747 (n_19473, n_4504, n_14265);
  nand g39748 (n_19458, n_4150, n_14202);
  nand g39749 (n_19470, n_4183, n_14233);
  nand g39750 (n_17709, n_14205, n_17708);
  nand g39751 (n_17714, \data_stack_mem[3] [5], n_11478);
  nand g39752 (n_17721, n_14224, n_17720);
  nand g39753 (n_4117, n_17660, n_17661);
  nand g39754 (n_19455, n_4471, n_14236);
  or g39755 (n_17661, wc404, n_14487);
  not gc404 (wc404, n_4085);
  nand g39756 (n_17720, \data_stack_mem[2] [6], n_12645);
  or g39757 (n_17660, n_4085, wc405);
  not gc405 (wc405, n_14487);
  nand g39758 (n_20780, n_14096, n_4151);
  or g39759 (n_20781, n_14096, n_4151);
  nand g39760 (n_4183, n_20780, n_20781);
  nand g39761 (n_17708, \data_stack_mem[4] [4], n_11540);
  nand g39762 (n_20782, n_14047, n_4184);
  or g39763 (n_20783, n_14047, n_4184);
  nand g39764 (n_4216, n_20782, n_20783);
  nand g39765 (n_11478, n_17615, n_19437);
  nand g39766 (n_17702, \data_stack_mem[5] [3], n_11673);
  nand g39767 (n_20784, n_14010, n_4118);
  or g39768 (n_20785, n_14010, n_4118);
  nand g39769 (n_4150, n_20784, n_20785);
  or g39770 (n_17647, \data_stack_mem[7] [1], wc406);
  not gc406 (wc406, n_13813);
  or g39771 (n_17648, wc407, n_13813);
  not gc407 (wc407, \data_stack_mem[7] [1]);
  or g39772 (n_17679, wc408, n_13791);
  not gc408 (wc408, data_stack_pointer[3]);
  nand g39773 (n_19446, n_4373, n_14222);
  nand g39774 (n_4372, n_17672, n_17673);
  or g39775 (n_17684, \data_stack_mem[2] [6], wc409);
  not gc409 (wc409, n_12722);
  or g39776 (n_17655, n_13400, wc410);
  not gc410 (wc410, n_13791);
  or g39777 (n_17654, n_13791, n_14151);
  or g39778 (n_17579, \data_stack_mem[4] [3], wc411);
  not gc411 (wc411, n_12166);
  nand g39779 (n_14491, n_17621, n_17622);
  nand g39780 (n_19422, n_4439, n_14208);
  or g39781 (n_17696, \data_stack_mem[6] [2], wc412);
  not gc412 (wc412, n_12317);
  nand g39782 (n_20786, n_14064, n_4472);
  or g39783 (n_20787, n_14064, n_4472);
  nand g39784 (n_4504, n_20786, n_20787);
  nand g39785 (n_17726, \data_stack_mem[6] [2], n_11723);
  or g39786 (n_17732, \data_stack_mem[7] [1], wc413);
  not gc413 (wc413, n_13791);
  nand g39787 (n_20788, n_14093, n_4439);
  or g39788 (n_20789, n_14093, n_4439);
  nand g39789 (n_4471, n_20788, n_20789);
  nand g39790 (n_4084, n_17666, n_17667);
  or g39791 (n_17672, wc414, n_4340);
  not gc414 (wc414, n_14509);
  nand g39792 (n_14487, n_17555, n_17556);
  or g39793 (n_17639, \data_stack_mem[3] [4], wc415);
  not gc415 (wc415, n_12045);
  nand g39794 (n_12645, n_17627, n_19440);
  nand g39795 (n_19437, n_4085, n_14221);
  nand g39796 (n_11723, n_17609, n_19434);
  or g39797 (n_17667, n_14504, wc416);
  not gc416 (wc416, n_4052);
  or g39798 (n_17666, wc417, n_4052);
  not gc417 (wc417, n_14504);
  nand g39799 (n_17678, n_14524, n_1409);
  nand g39800 (n_12722, n_17633, n_19443);
  or g39801 (n_17622, n_13766, wc418);
  not gc418 (wc418, n_12045);
  or g39802 (n_17621, n_14133, n_12045);
  or g39803 (n_14047, n_17610, n_3910);
  or g39804 (n_14010, n_20, n_17604);
  nand g39805 (n_20790, n_14029, n_4407);
  or g39806 (n_20791, n_14029, n_4407);
  nand g39807 (n_4439, n_20790, n_20791);
  or g39808 (n_14093, n_17586, n_3908);
  nand g39809 (n_11540, n_17603, n_19431);
  nand g39810 (n_12317, n_17591, n_19425);
  nand g39811 (n_11673, n_17597, n_19428);
  or g39812 (n_14064, n_17592, n_3910);
  nand g39813 (n_20792, n_14053, n_4374);
  or g39814 (n_20793, n_14053, n_4374);
  nand g39815 (n_4406, n_20792, n_20793);
  or g39816 (n_14096, n_17598, n_3908);
  or g39817 (n_17673, n_14509, wc419);
  not gc419 (wc419, n_4340);
  nand g39818 (n_12166, n_17507, n_19395);
  nand g39819 (n_19428, n_4151, n_14206);
  nand g39820 (n_19434, n_4184, n_14199);
  nand g39821 (n_17592, n_14200, n_17591);
  nand g39822 (n_17604, n_14212, n_17603);
  nand g39823 (n_19431, n_4118, n_14212);
  nand g39824 (n_17586, n_14208, n_17585);
  nand g39825 (n_19425, n_4472, n_14200);
  or g39826 (n_17555, n_13766, n_11449);
  or g39827 (n_17556, n_14133, wc420);
  not gc420 (wc420, n_11449);
  nand g39828 (n_17615, \data_stack_mem[3] [4], n_11449);
  nand g39829 (n_19395, n_14223, n_4407);
  nand g39830 (n_14504, n_17561, n_17562);
  nand g39831 (n_19440, n_14231, n_4052);
  nand g39832 (n_17598, n_14206, n_17597);
  nand g39833 (n_1409, n_17573, n_17574);
  or g39834 (n_14029, n_20, n_17508);
  nand g39835 (n_17610, n_14199, n_17609);
  nand g39836 (n_12045, n_17549, n_19416);
  nand g39837 (n_14509, n_17567, n_17568);
  or g39838 (n_14053, wc421, n_17550);
  not gc421 (wc421, n_37);
  nand g39839 (n_19443, n_14273, n_4340);
  nand g39840 (n_20794, n_14049, n_4119);
  or g39841 (n_20795, n_14049, n_4119);
  nand g39842 (n_4151, n_20794, n_20795);
  nand g39843 (n_17597, \data_stack_mem[5] [2], n_11622);
  nand g39844 (n_20796, n_14072, n_4440);
  or g39845 (n_20797, n_14072, n_4440);
  nand g39846 (n_4472, n_20796, n_20797);
  or g39847 (n_4407, wc422, n_17478);
  not gc422 (wc422, n_17477);
  or g39848 (n_17633, \data_stack_mem[2] [5], wc423);
  not gc423 (wc423, n_12720);
  nand g39849 (n_17550, n_14227, n_17549);
  or g39850 (n_17568, n_13912, wc424);
  not gc424 (wc424, n_12720);
  or g39851 (n_17567, n_13821, n_12720);
  nand g39852 (n_20798, n_14056, n_4341);
  or g39853 (n_20799, n_14056, n_4341);
  nand g39854 (n_4373, n_20798, n_20799);
  nand g39855 (n_11449, n_17537, n_19410);
  nand g39856 (n_19416, n_14227, n_4374);
  nand g39857 (n_20800, n_14051, n_4053);
  or g39858 (n_20801, n_14051, n_4053);
  nand g39859 (n_4085, n_20800, n_20801);
  or g39860 (n_17609, wc425, n_13807);
  not gc425 (wc425, \data_stack_mem[6] [1]);
  or g39861 (n_17585, \data_stack_mem[5] [2], wc426);
  not gc426 (wc426, n_12218);
  nand g39862 (n_17508, n_14223, n_17507);
  or g39863 (n_17574, n_13783, n_3910);
  nand g39864 (n_20802, n_14052, n_4086);
  or g39865 (n_20803, n_14052, n_4086);
  nand g39866 (n_4118, n_20802, n_20803);
  nand g39867 (n_17627, \data_stack_mem[2] [5], n_12643);
  or g39868 (n_17591, \data_stack_mem[6] [1], wc427);
  not gc427 (wc427, n_13783);
  or g39869 (n_17562, n_13821, wc428);
  not gc428 (wc428, n_12643);
  or g39870 (n_17561, n_13912, n_12643);
  nand g39871 (n_20804, n_14034, n_4152);
  or g39872 (n_20805, n_14034, n_4152);
  nand g39873 (n_4184, n_20804, n_20805);
  nand g39874 (n_17603, \data_stack_mem[4] [3], n_11572);
  nand g39875 (n_17477, n_14466, n_4375);
  or g39876 (n_17507, \data_stack_mem[4] [2], wc429);
  not gc429 (wc429, n_12119);
  nand g39877 (n_12720, n_17513, n_19398);
  or g39878 (n_14056, n_17514, wc430);
  not gc430 (wc430, n_3902);
  nand g39879 (n_12218, n_17519, n_19401);
  or g39880 (n_17549, \data_stack_mem[3] [3], wc431);
  not gc431 (wc431, n_12070);
  or g39881 (n_14034, n_17526, n_3908);
  nand g39882 (n_17573, n_14196, n_1393);
  or g39883 (n_14049, n_20, n_17532);
  nand g39884 (n_12643, n_17543, n_19413);
  or g39885 (n_14072, n_17520, n_3908);
  nand g39886 (n_19410, n_14292, n_4086);
  or g39887 (n_14051, n_17544, wc432);
  not gc432 (wc432, n_3902);
  or g39888 (n_14052, wc433, n_17538);
  not gc433 (wc433, n_37);
  nand g39889 (n_11622, n_17525, n_19404);
  nand g39890 (n_11572, n_17531, n_19407);
  nand g39891 (n_17478, n_17475, n_17476);
  nand g39892 (n_12070, n_17495, n_17496);
  nand g39893 (n_17514, n_14249, n_17513);
  nand g39894 (n_19413, n_4053, n_14258);
  nand g39895 (n_1393, n_17501, n_17502);
  nand g39896 (n_19401, n_4440, n_14216);
  nand g39897 (n_17544, n_14258, n_17543);
  nand g39898 (n_17532, n_14220, n_17531);
  nand g39899 (n_17526, n_14215, n_17525);
  nand g39900 (n_17520, n_14216, n_17519);
  or g39901 (n_14466, wc434, n_17385);
  not gc434 (wc434, n_37);
  nand g39902 (n_12119, n_17423, n_19383);
  nand g39903 (n_17538, n_14292, n_17537);
  nand g39904 (n_19404, n_4152, n_14215);
  or g39905 (n_4086, wc435, n_17457);
  not gc435 (wc435, n_17456);
  nand g39906 (n_19398, n_4341, n_14249);
  nand g39907 (n_19407, n_14220, n_4119);
  or g39908 (n_17502, n_3908, n_13781);
  nand g39909 (n_20806, n_14069, n_4408);
  or g39910 (n_20807, n_14069, n_4408);
  nand g39911 (n_4440, n_20806, n_20807);
  nand g39912 (n_20808, n_14041, n_4120);
  or g39913 (n_20809, n_14041, n_4120);
  nand g39914 (n_4152, n_20808, n_20809);
  or g39915 (n_17519, \data_stack_mem[5] [1], wc436);
  not gc436 (wc436, n_13781);
  nand g39916 (n_17531, \data_stack_mem[4] [2], n_11521);
  or g39917 (n_17475, n_14130, n_14288);
  nand g39918 (n_17385, n_17383, n_17384);
  nand g39919 (n_19383, n_14270, n_4408);
  nand g39920 (n_4330, n_14578, n_3793);
  or g39921 (n_17513, \data_stack_mem[2] [4], wc437);
  not gc437 (wc437, n_12699);
  nand g39922 (n_4119, n_17483, n_17484);
  nand g39923 (n_4374, n_17489, n_17490);
  or g39924 (n_17495, \data_stack_mem[3] [2], wc438);
  not gc438 (wc438, n_14288);
  or g39925 (n_17525, wc439, n_13805);
  not gc439 (wc439, \data_stack_mem[5] [1]);
  or g39926 (n_4050, wc440, n_15975);
  not gc440 (wc440, n_13987);
  nand g39927 (n_17543, \data_stack_mem[2] [4], n_12622);
  nand g39928 (n_17456, n_14485, n_4054);
  nand g39929 (n_17537, \data_stack_mem[3] [3], n_11474);
  or g39930 (n_4338, wc441, n_15984);
  not gc441 (wc441, n_13987);
  nand g39931 (n_11474, n_17435, n_19389);
  or g39932 (n_17384, wc442, n_12027);
  not gc442 (wc442, \data_stack_mem[3] [2]);
  nand g39933 (n_11521, n_17429, n_19386);
  or g39934 (n_17489, wc443, n_4342);
  not gc443 (wc443, n_14499);
  or g39935 (n_4051, wc444, n_15591);
  not gc444 (wc444, n_14134);
  or g39936 (n_14041, n_20, n_17430);
  or g39937 (n_17490, n_14499, wc445);
  not gc445 (wc445, n_4342);
  nand g39938 (n_14578, n_14673, n_19353);
  nand g39939 (n_15975, n_15973, n_15974);
  or g39940 (n_14485, n_17400, wc446);
  not gc446 (wc446, n_3902);
  or g39941 (n_4408, wc447, n_17370);
  not gc447 (wc447, n_17369);
  or g39942 (n_4339, wc448, n_15579);
  not gc448 (wc448, n_14134);
  or g39943 (n_14069, n_20, n_17424);
  nand g39944 (n_4049, n_19361, n_19362);
  nand g39945 (n_12699, n_17441, n_19392);
  nand g39946 (n_17501, n_14209, n_1377);
  nand g39947 (n_17457, n_17454, n_17455);
  nand g39948 (n_17496, n_4375, n_12027);
  or g39949 (n_17484, wc449, n_14479);
  not gc449 (wc449, n_4087);
  or g39950 (n_17476, n_17474, wc450);
  not gc450 (wc450, n_12027);
  or g39951 (n_17383, \data_stack_mem[3] [2], wc451);
  not gc451 (wc451, n_12027);
  nand g39952 (n_12622, n_17462, n_17463);
  nand g39953 (n_15984, n_15982, n_15983);
  or g39954 (n_17483, n_4087, wc452);
  not gc452 (wc452, n_14479);
  nand g39955 (n_17430, n_14263, n_17429);
  or g39956 (n_5685, n_17201, n_17202);
  nand g39957 (n_19389, n_4087, n_14234);
  or g39958 (n_5669, n_16769, n_16770);
  or g39959 (n_5683, n_16337, n_16338);
  or g39960 (n_5711, n_16721, n_16722);
  or g39961 (n_5687, n_17153, n_17154);
  or g39962 (n_5661, n_17249, n_17250);
  or g39963 (n_5681, n_16385, n_16386);
  or g39964 (n_5689, n_17105, n_17106);
  nand g39965 (n_17400, n_17398, n_17399);
  or g39966 (n_5673, n_17057, n_17058);
  or g39967 (n_5667, n_16817, n_16818);
  nand g39968 (n_19386, n_4120, n_14263);
  nand g39969 (n_12027, n_17375, n_17376);
  or g39970 (n_5663, n_17297, n_17298);
  nand g39971 (n_14499, n_17405, n_17406);
  or g39972 (n_17454, n_13803, n_14269);
  or g39973 (n_5679, n_16433, n_16434);
  nand g39974 (n_17424, n_14270, n_17423);
  or g39975 (n_5695, n_16673, n_16674);
  or g39976 (n_5657, n_16961, n_16962);
  nand g39977 (n_19392, n_14284, n_4342);
  or g39978 (n_5677, n_16481, n_16482);
  nand g39979 (n_1377, n_17417, n_17418);
  or g39980 (n_5665, n_16865, n_16866);
  or g39981 (n_5655, n_17009, n_17010);
  or g39982 (n_5659, n_16913, n_16914);
  or g39983 (n_5709, n_16625, n_16626);
  or g39984 (n_19362, n_14173, wc453);
  not gc453 (wc453, n_14567);
  or g39985 (n_17474, n_4375, n_13767);
  nand g39986 (n_15579, n_15577, n_15578);
  or g39987 (n_5693, n_16577, n_16578);
  or g39988 (n_15974, wc454, n_14192);
  not gc454 (wc454, n_14567);
  nand g39989 (n_14479, n_17390, n_17391);
  nand g39990 (n_17370, n_17367, n_17368);
  or g39991 (n_15973, n_13898, n_14567);
  nand g39992 (n_15591, n_15589, n_15590);
  or g39993 (n_5675, n_16529, n_16530);
  or g39994 (n_15982, n_13898, n_14572);
  or g39995 (n_15983, wc455, n_14192);
  not gc455 (wc455, n_14572);
  nand g39996 (n_19353, n_14572, n_14170);
  nand g39997 (n_17462, \data_stack_mem[2] [3], n_14269);
  or g39998 (n_16962, n_16959, n_16960);
  or g39999 (n_17423, \data_stack_mem[4] [1], wc456);
  not gc456 (wc456, n_13779);
  nand g40000 (n_14572, n_13935, n_15600);
  or g40001 (n_15589, n_15588, wc457);
  not gc457 (wc457, n_3793);
  or g40002 (n_16578, n_16575, n_16576);
  nand g40003 (n_17369, n_14475, n_4376);
  or g40004 (n_17010, n_17007, n_17008);
  nand g40005 (n_14567, n_13938, n_15597);
  or g40006 (n_17367, n_17366, wc458);
  not gc458 (wc458, n_13788);
  or g40007 (n_17368, n_14153, n_14242);
  or g40008 (n_16530, n_16527, n_16528);
  or g40009 (n_17391, n_14130, wc459);
  not gc459 (wc459, n_11432);
  or g40010 (n_15578, n_15576, wc460);
  not gc460 (wc460, n_3793);
  or g40011 (n_17390, n_13767, n_11432);
  or g40012 (n_16626, n_16623, n_16624);
  or g40013 (n_16914, n_16911, n_16912);
  or g40014 (n_17418, n_20, n_13779);
  or g40015 (n_16866, n_16863, n_16864);
  or g40016 (n_16482, n_16479, n_16480);
  or g40017 (n_16674, n_16671, n_16672);
  or g40018 (n_17441, \data_stack_mem[2] [3], wc461);
  not gc461 (wc461, n_12716);
  nand g40019 (n_17463, n_4054, n_12639);
  or g40020 (n_17455, n_17453, wc462);
  not gc462 (wc462, n_12639);
  or g40021 (n_17406, n_13803, wc463);
  not gc463 (wc463, n_12716);
  or g40022 (n_17405, n_14126, n_12716);
  or g40023 (n_16434, n_16431, n_16432);
  or g40024 (n_17298, n_17295, n_17296);
  nand g40025 (n_17435, \data_stack_mem[3] [2], n_11432);
  or g40026 (n_17375, \data_stack_mem[3] [1], wc464);
  not gc464 (wc464, n_14242);
  nand g40027 (n_20810, n_14054, n_4343);
  or g40028 (n_20811, n_14054, n_4343);
  nand g40029 (n_4375, n_20810, n_20811);
  or g40030 (n_17058, n_17055, n_17056);
  nand g40031 (n_20812, n_14076, n_4055);
  or g40032 (n_20813, n_14076, n_4055);
  nand g40033 (n_4087, n_20812, n_20813);
  or g40034 (n_17106, n_17103, n_17104);
  nand g40035 (n_4120, n_17411, n_17412);
  nand g40036 (n_17399, \data_stack_mem[2] [3], n_12639);
  or g40037 (n_17398, \data_stack_mem[2] [3], n_12639);
  or g40038 (n_16386, n_16383, n_16384);
  or g40039 (n_17250, n_17247, n_17248);
  or g40040 (n_17154, n_17151, n_17152);
  or g40041 (n_16818, n_16815, n_16816);
  or g40042 (n_16722, n_16719, n_16720);
  or g40043 (n_16338, n_16335, n_16336);
  or g40044 (n_17202, n_17199, n_17200);
  or g40045 (n_5653, n_16265, n_16266);
  or g40046 (n_16770, n_16767, n_16768);
  or g40047 (n_17429, wc465, n_13798);
  not gc465 (wc465, \data_stack_mem[4] [1]);
  or g40048 (n_15577, n_14144, n_13123);
  nand g40049 (n_4880, n_16007, n_16008);
  or g40050 (n_16336, wc466, n_16332);
  not gc466 (wc466, n_16331);
  or g40051 (n_17201, n_17197, n_17198);
  or g40052 (n_17200, wc467, n_17196);
  not gc467 (wc467, n_17195);
  or g40053 (n_16337, n_16333, n_16334);
  or g40054 (n_18671, n_18667, wc468);
  not gc468 (wc468, \data_stack_mem[8] [5]);
  nand g40055 (n_15576, n_1326, n_13123);
  nand g40056 (n_4768, n_16163, n_16164);
  or g40057 (n_16266, n_16263, n_16264);
  or g40058 (n_16720, wc469, n_16716);
  not gc469 (wc469, n_16715);
  or g40059 (n_16672, wc470, n_16668);
  not gc470 (wc470, n_16667);
  or g40060 (n_16265, n_16261, n_16262);
  nand g40061 (n_4828, n_15713, n_15714);
  nand g40062 (n_4804, n_16187, n_16188);
  or g40063 (n_17248, wc471, n_17244);
  not gc471 (wc471, n_17243);
  nand g40064 (n_4876, n_16001, n_16002);
  or g40065 (n_17153, n_17149, n_17150);
  nand g40066 (n_4904, n_16043, n_16044);
  nand g40067 (n_11432, n_17315, n_19380);
  or g40068 (n_17152, wc472, n_17148);
  not gc472 (wc472, n_17147);
  nand g40069 (n_4844, n_15845, n_15846);
  or g40070 (n_16673, n_16669, n_16670);
  or g40071 (n_16384, wc473, n_16380);
  not gc473 (wc473, n_16379);
  or g40072 (n_16385, n_16381, n_16382);
  or g40073 (n_18782, n_18778, wc474);
  not gc474 (wc474, \data_stack_mem[8] [6]);
  nand g40074 (n_4752, n_16139, n_16140);
  or g40075 (n_17249, n_17245, n_17246);
  or g40076 (n_17009, n_17005, n_17006);
  or g40077 (n_17008, wc475, n_17004);
  not gc475 (wc475, n_17003);
  nand g40078 (n_15597, n_13774, n_11318);
  or g40079 (n_17412, n_14482, wc476);
  not gc476 (wc476, n_4088);
  nand g40080 (n_4796, n_16223, n_16224);
  or g40081 (n_17105, n_17101, n_17102);
  or g40082 (n_17104, wc477, n_17100);
  not gc477 (wc477, n_17099);
  nand g40083 (n_4900, n_16037, n_16038);
  or g40084 (n_16817, n_16813, n_16814);
  or g40085 (n_3711, n_3710, wc478);
  not gc478 (wc478, n_14589);
  or g40086 (n_16816, wc479, n_16812);
  not gc479 (wc479, n_16811);
  or g40087 (n_15600, wc480, n_13123);
  not gc480 (wc480, n_13780);
  nand g40088 (n_4896, n_16031, n_16032);
  or g40089 (n_16721, n_16717, n_16718);
  or g40090 (n_16576, wc481, n_16572);
  not gc481 (wc481, n_16571);
  or g40091 (n_17057, n_17053, n_17054);
  or g40092 (n_17056, wc482, n_17052);
  not gc482 (wc482, n_17051);
  or g40093 (n_15590, n_14144, wc483);
  not gc483 (wc483, n_11318);
  or g40094 (n_15588, wc484, n_11318);
  not gc484 (wc484, n_1326);
  or g40095 (n_16624, wc485, n_16620);
  not gc485 (wc485, n_16619);
  nand g40096 (n_4892, n_16025, n_16026);
  or g40097 (n_16432, wc486, n_16428);
  not gc486 (wc486, n_16427);
  or g40098 (n_16865, n_16861, n_16862);
  or g40099 (n_14054, n_16284, wc487);
  not gc487 (wc487, n_3902);
  or g40100 (n_16625, n_16621, n_16622);
  or g40101 (n_16433, n_16429, n_16430);
  or g40102 (n_16864, wc488, n_16860);
  not gc488 (wc488, n_16859);
  nand g40103 (n_4800, n_16217, n_16218);
  nand g40104 (n_17376, n_13788, n_4376);
  or g40105 (n_17296, wc489, n_17292);
  not gc489 (wc489, n_17291);
  nand g40106 (n_4816, n_15701, n_15702);
  or g40107 (n_17297, n_17293, n_17294);
  or g40108 (n_16768, wc490, n_16764);
  not gc490 (wc490, n_16763);
  nand g40109 (n_4764, n_16157, n_16158);
  nand g40110 (n_12716, n_16283, n_19374);
  nand g40111 (n_4848, n_15851, n_15852);
  nand g40112 (n_4780, n_16211, n_16212);
  or g40113 (n_16961, n_16957, n_16958);
  nand g40114 (n_4748, n_16133, n_16134);
  nand g40115 (n_4840, n_15719, n_15720);
  nand g40116 (n_4784, n_16205, n_16206);
  nand g40117 (n_12639, n_16289, n_19377);
  nand g40118 (n_4852, n_15857, n_15858);
  nand g40119 (n_4788, n_16199, n_16200);
  or g40120 (n_16960, wc491, n_16956);
  not gc491 (wc491, n_16955);
  nand g40121 (n_4756, n_16145, n_16146);
  nand g40122 (n_4856, n_15863, n_15864);
  nand g40123 (n_4808, n_16181, n_16182);
  nand g40124 (n_4812, n_15725, n_15726);
  or g40125 (n_16913, n_16909, n_16910);
  nand g40126 (n_4860, n_15869, n_15870);
  or g40127 (n_16480, wc492, n_16476);
  not gc492 (wc492, n_16475);
  or g40128 (n_4052, wc493, n_15465);
  not gc493 (wc493, n_14160);
  nand g40129 (n_4868, n_15881, n_15882);
  nand g40130 (n_17417, n_14226, n_1361);
  nand g40131 (n_4864, n_15875, n_15876);
  nand g40132 (n_4824, n_15731, n_15732);
  or g40133 (n_16577, n_16573, n_16574);
  or g40134 (n_3684, wc494, n_3683);
  not gc494 (wc494, n_14591);
  nand g40135 (n_4792, n_16193, n_16194);
  nand g40136 (n_4820, n_15707, n_15708);
  or g40137 (n_16912, wc495, n_16908);
  not gc495 (wc495, n_16907);
  or g40138 (n_17411, wc496, n_4088);
  not gc496 (wc496, n_14482);
  nand g40139 (n_4872, n_15887, n_15888);
  or g40140 (n_16528, wc497, n_16524);
  not gc497 (wc497, n_16523);
  or g40141 (n_16481, n_16477, n_16478);
  or g40142 (n_14475, wc498, n_15945);
  not gc498 (wc498, n_37);
  or g40143 (n_18123, n_18121, wc499);
  not gc499 (wc499, \data_stack_mem[8] [1]);
  nand g40144 (n_4760, n_16151, n_16152);
  or g40145 (n_16529, n_16525, n_16526);
  or g40146 (n_17366, n_4376, n_13764);
  or g40147 (n_4340, wc500, n_15474);
  not gc500 (wc500, n_14160);
  nand g40148 (n_4776, n_16175, n_16176);
  or g40149 (n_14076, n_16290, wc501);
  not gc501 (wc501, n_3902);
  nand g40150 (n_4888, n_16019, n_16020);
  or g40151 (n_17858, n_3673, wc502);
  not gc502 (wc502, n_14240);
  nand g40152 (n_4832, n_15737, n_15738);
  nand g40153 (n_4772, n_16169, n_16170);
  nand g40154 (n_4884, n_16013, n_16014);
  or g40155 (n_18428, n_18424, wc503);
  not gc503 (wc503, \data_stack_mem[8] [3]);
  nand g40156 (n_4836, n_15743, n_15744);
  or g40157 (n_16769, n_16765, n_16766);
  nand g40158 (n_16764, n_16755, n_16756);
  nand g40159 (n_16332, n_16323, n_16324);
  nand g40160 (n_17198, n_17191, n_17192);
  nand g40161 (n_17244, n_17235, n_17236);
  nand g40162 (n_17196, n_17187, n_17188);
  nand g40163 (n_17246, n_17239, n_17240);
  nand g40164 (n_16380, n_16371, n_16372);
  nand g40165 (n_16382, n_16375, n_16376);
  nand g40166 (n_4744, n_15791, n_15792);
  nand g40167 (n_4968, n_15797, n_15798);
  nand g40168 (n_16044, \data_stack_mem[6] [7], n_13111);
  nand g40169 (n_4956, n_15803, n_15804);
  nand g40170 (n_4960, n_15809, n_15810);
  nand g40171 (n_17150, n_17143, n_17144);
  nand g40172 (n_17148, n_17139, n_17140);
  nand g40173 (n_16263, n_16257, n_16258);
  nand g40174 (n_16428, n_16419, n_16420);
  nand g40175 (n_16261, n_16253, n_16254);
  nand g40176 (n_17102, n_17095, n_17096);
  nand g40177 (n_16038, \data_stack_mem[6] [6], n_13111);
  nand g40178 (n_17100, n_17091, n_17092);
  nand g40179 (n_16430, n_16423, n_16424);
  nand g40180 (n_17292, n_17283, n_17284);
  nand g40181 (n_16224, \data_stack_mem[3] [4], n_13110);
  nand g40182 (n_16032, \data_stack_mem[6] [5], n_13111);
  nand g40183 (n_16140, \data_stack_mem[2] [1], n_13106);
  nand g40184 (n_17054, n_17047, n_17048);
  nand g40185 (n_16284, n_14244, n_16283);
  nand g40186 (n_17294, n_17287, n_17288);
  or g40187 (n_4376, wc504, n_15621);
  not gc504 (wc504, n_15620);
  nand g40188 (n_4928, n_15659, n_15660);
  nand g40189 (n_15720, \data_stack_mem[4] [7], n_13108);
  nand g40190 (n_19374, n_4343, n_14244);
  nand g40191 (n_16218, \data_stack_mem[3] [5], n_13110);
  nand g40192 (n_16212, \data_stack_mem[3] [0], n_13110);
  or g40193 (n_18315, n_18313, wc505);
  not gc505 (wc505, \data_stack_mem[8] [2]);
  nand g40194 (n_16206, \data_stack_mem[3] [1], n_13110);
  nand g40195 (n_4924, n_15653, n_15654);
  nand g40196 (n_15726, \data_stack_mem[4] [0], n_13108);
  nand g40197 (n_16476, n_16467, n_16468);
  or g40198 (n_4341, wc506, n_15276);
  not gc506 (wc506, n_13981);
  nand g40199 (n_16478, n_16471, n_16472);
  nand g40200 (n_17052, n_17043, n_17044);
  nand g40201 (n_16766, n_16759, n_16760);
  nand g40202 (n_1361, n_15989, n_15990);
  nand g40203 (n_15732, \data_stack_mem[4] [3], n_13108);
  nand g40204 (n_16200, \data_stack_mem[3] [2], n_13110);
  nand g40205 (n_15714, \data_stack_mem[4] [4], n_13108);
  nand g40206 (n_16524, n_16515, n_16516);
  nand g40207 (n_4952, n_15815, n_15816);
  nand g40208 (n_16526, n_16519, n_16520);
  nand g40209 (n_4948, n_15821, n_15822);
  nand g40210 (n_15474, n_15472, n_15473);
  or g40211 (n_18121, n_1427, n_13900);
  nand g40212 (n_4944, n_15827, n_15828);
  nand g40213 (n_18126, n_14553, n_1427);
  nand g40214 (n_16026, \data_stack_mem[6] [4], n_13111);
  nand g40215 (n_15738, \data_stack_mem[4] [5], n_13108);
  nand g40216 (n_16020, \data_stack_mem[6] [3], n_13111);
  nand g40217 (n_15708, \data_stack_mem[4] [2], n_13108);
  nand g40218 (n_16014, \data_stack_mem[6] [2], n_13111);
  nand g40219 (n_13123, n_14670, n_19350);
  nand g40220 (n_4940, n_15833, n_15834);
  nand g40221 (n_16008, \data_stack_mem[6] [1], n_13111);
  nand g40222 (n_4964, n_15839, n_15840);
  nand g40223 (n_16194, \data_stack_mem[3] [3], n_13110);
  nand g40224 (n_15846, \data_stack_mem[5] [0], n_13107);
  or g40225 (n_14551, n_3673, wc507);
  not gc507 (wc507, n_15135);
  nand g40226 (n_14482, n_15950, n_15951);
  nand g40227 (n_17006, n_16999, n_17000);
  nand g40228 (n_16572, n_16563, n_16564);
  nand g40229 (n_17004, n_16995, n_16996);
  nand g40230 (n_16574, n_16567, n_16568);
  or g40231 (n_14552, n_12739, n_15372);
  nand g40232 (n_11318, n_14925, n_19368);
  nand g40233 (n_16002, \data_stack_mem[6] [0], n_13111);
  nand g40234 (n_16188, \data_stack_mem[3] [6], n_13110);
  nand g40235 (n_16134, \data_stack_mem[2] [0], n_13106);
  nand g40236 (n_15702, \data_stack_mem[4] [1], n_13108);
  nand g40237 (n_15852, \data_stack_mem[5] [1], n_13107);
  nand g40238 (n_15858, \data_stack_mem[5] [2], n_13107);
  nand g40239 (n_15864, \data_stack_mem[5] [3], n_13107);
  nand g40240 (n_15870, \data_stack_mem[5] [4], n_13107);
  nand g40241 (n_15876, \data_stack_mem[5] [5], n_13107);
  nand g40242 (n_3683, n_15446, n_15447);
  or g40243 (n_19041, n_19039, wc508);
  not gc508 (wc508, \data_stack_mem[8] [7]);
  nand g40244 (n_15465, n_15463, n_15464);
  nand g40245 (n_15945, n_15943, n_15944);
  nand g40246 (n_16182, \data_stack_mem[3] [7], n_13110);
  nand g40247 (n_16176, \data_stack_mem[2] [7], n_13106);
  nand g40248 (n_4916, n_15695, n_15696);
  nand g40249 (n_15744, \data_stack_mem[4] [6], n_13108);
  nand g40250 (n_16170, \data_stack_mem[2] [6], n_13106);
  nand g40251 (n_4920, n_15689, n_15690);
  nand g40252 (n_16164, \data_stack_mem[2] [5], n_13106);
  nand g40253 (n_18783, n_14495, n_1437);
  nand g40254 (n_15882, \data_stack_mem[5] [6], n_13107);
  or g40255 (n_18778, n_1437, n_13900);
  nand g40256 (n_16620, n_16611, n_16612);
  nand g40257 (n_19380, n_4088, n_14243);
  nand g40258 (n_16622, n_16615, n_16616);
  nand g40259 (n_4716, n_15749, n_15750);
  nand g40260 (n_16958, n_16951, n_16952);
  nand g40261 (n_16956, n_16947, n_16948);
  nand g40262 (n_4908, n_15683, n_15684);
  nand g40263 (n_16290, n_14289, n_16289);
  or g40264 (n_4053, wc509, n_15264);
  not gc509 (wc509, n_13981);
  nand g40265 (n_15888, \data_stack_mem[5] [7], n_13107);
  nand g40266 (n_16668, n_16659, n_16660);
  nand g40267 (n_16910, n_16903, n_16904);
  nand g40268 (n_16670, n_16663, n_16664);
  or g40269 (n_18667, n_1435, n_13900);
  nand g40270 (n_4696, n_15893, n_15894);
  nand g40271 (n_16908, n_16899, n_16900);
  nand g40272 (n_4692, n_15899, n_15900);
  nand g40273 (n_4684, n_15905, n_15906);
  nand g40274 (n_18672, n_14512, n_1435);
  nand g40275 (n_16158, \data_stack_mem[2] [4], n_13106);
  nand g40276 (n_4932, n_15677, n_15678);
  nand g40277 (n_4936, n_15665, n_15666);
  nand g40278 (n_16862, n_16855, n_16856);
  nand g40279 (n_16146, \data_stack_mem[2] [2], n_13106);
  nand g40280 (n_16860, n_16851, n_16852);
  or g40281 (n_14240, n_15021, wc510);
  not gc510 (wc510, n_14226);
  or g40282 (n_3693, wc511, n_3692);
  not gc511 (wc511, n_14586);
  nand g40283 (n_3710, n_15440, n_15441);
  nand g40284 (n_4700, n_15935, n_15936);
  nand g40285 (n_4720, n_15755, n_15756);
  nand g40286 (n_4740, n_15785, n_15786);
  nand g40287 (n_16152, \data_stack_mem[2] [3], n_13106);
  nand g40288 (n_4724, n_15761, n_15762);
  nand g40289 (n_4704, n_15929, n_15930);
  nand g40290 (n_18429, n_14532, n_1431);
  nand g40291 (n_16716, n_16707, n_16708);
  nand g40292 (n_16718, n_16711, n_16712);
  or g40293 (n_18424, n_1431, n_13900);
  nand g40294 (n_16814, n_16807, n_16808);
  nand g40295 (n_16812, n_16803, n_16804);
  nand g40296 (n_19377, n_4055, n_14289);
  nand g40297 (n_4736, n_15779, n_15780);
  nand g40298 (n_4912, n_15671, n_15672);
  nand g40299 (n_4688, n_15911, n_15912);
  nand g40300 (n_4732, n_15773, n_15774);
  nand g40301 (n_4708, n_15917, n_15918);
  nand g40302 (n_4728, n_15767, n_15768);
  nand g40303 (n_4712, n_15923, n_15924);
  nand g40304 (n_16334, n_16327, n_16328);
  nand g40305 (n_3692, n_15434, n_15435);
  nand g40306 (n_16765, n_16757, n_16758);
  nand g40307 (n_15930, \data_stack_mem[0] [5], n_13109);
  or g40308 (n_16760, wc512, n_13405);
  not gc512 (wc512, \out_fifo[4][0] [8]);
  nand g40309 (n_15767, \data_stack_mem[1] [3], n_12808);
  nand g40310 (n_16767, n_16761, n_16762);
  nand g40311 (n_15773, \data_stack_mem[1] [4], n_12808);
  nand g40312 (n_15924, \data_stack_mem[0] [7], n_13109);
  nand g40313 (n_15779, \data_stack_mem[1] [5], n_12808);
  nand g40314 (n_15918, \data_stack_mem[0] [6], n_13109);
  or g40315 (n_16756, wc513, n_13770);
  not gc513 (wc513, \out_fifo[0][0] [8]);
  or g40316 (n_16804, wc514, n_13770);
  not gc514 (wc514, \out_fifo[0][0] [7]);
  or g40317 (n_16808, wc515, n_13405);
  not gc515 (wc515, \out_fifo[4][0] [7]);
  nand g40318 (n_16813, n_16805, n_16806);
  nand g40319 (n_16815, n_16809, n_16810);
  nand g40320 (n_16719, n_16713, n_16714);
  nand g40321 (n_20814, n_13965, n_1415);
  or g40322 (n_20815, n_13965, n_1415);
  nand g40323 (n_1431, n_20814, n_20815);
  nand g40324 (n_16717, n_16709, n_16710);
  nand g40325 (n_15785, \data_stack_mem[1] [6], n_12808);
  nand g40326 (n_15912, \data_stack_mem[0] [1], n_13109);
  or g40327 (n_16712, wc516, n_13405);
  not gc516 (wc516, \out_fifo[4][2] [9]);
  or g40328 (n_16708, wc517, n_13770);
  not gc517 (wc517, \out_fifo[0][2] [9]);
  or g40329 (n_16852, wc518, n_13770);
  not gc518 (wc518, \out_fifo[0][0] [6]);
  or g40330 (n_16856, wc519, n_13405);
  not gc519 (wc519, \out_fifo[4][0] [6]);
  nand g40331 (n_15936, \data_stack_mem[0] [4], n_13109);
  nand g40332 (n_15761, \data_stack_mem[1] [2], n_12808);
  or g40333 (n_15440, wc520, n_3673);
  not gc520 (wc520, n_14588);
  nand g40334 (n_16861, n_16853, n_16854);
  nand g40335 (n_16863, n_16857, n_16858);
  or g40336 (n_16900, wc521, n_13770);
  not gc521 (wc521, \out_fifo[0][0] [3]);
  nand g40337 (n_15906, \data_stack_mem[0] [0], n_13109);
  nand g40338 (n_16671, n_16665, n_16666);
  or g40339 (n_16904, wc522, n_13405);
  not gc522 (wc522, \out_fifo[4][0] [3]);
  nand g40340 (n_15900, \data_stack_mem[0] [2], n_13109);
  nand g40341 (n_20816, n_13958, n_1419);
  or g40342 (n_20817, n_13958, n_1419);
  nand g40343 (n_1435, n_20816, n_20817);
  nand g40344 (n_15894, \data_stack_mem[0] [3], n_13109);
  nand g40345 (n_16669, n_16661, n_16662);
  nand g40346 (n_16909, n_16901, n_16902);
  or g40347 (n_16664, wc523, n_13405);
  not gc523 (wc523, \out_fifo[4][2] [1]);
  or g40348 (n_16660, wc524, n_13770);
  not gc524 (wc524, \out_fifo[0][2] [1]);
  nand g40349 (n_16911, n_16905, n_16906);
  or g40350 (n_16948, wc525, n_13770);
  not gc525 (wc525, \out_fifo[0][0] [2]);
  or g40351 (n_16952, wc526, n_13405);
  not gc526 (wc526, \out_fifo[4][0] [2]);
  nand g40352 (n_16957, n_16949, n_16950);
  nand g40353 (n_16623, n_16617, n_16618);
  nand g40354 (n_15755, \data_stack_mem[1] [1], n_12808);
  nand g40355 (n_5787, n_16097, n_16098);
  nand g40356 (n_16621, n_16613, n_16614);
  nand g40357 (n_16959, n_16953, n_16954);
  or g40358 (n_16616, wc527, n_13405);
  not gc527 (wc527, \out_fifo[4][2] [8]);
  or g40359 (n_16612, wc528, n_13770);
  not gc528 (wc528, \out_fifo[0][2] [8]);
  nand g40360 (n_20818, n_13959, n_1421);
  or g40361 (n_20819, n_13959, n_1421);
  nand g40362 (n_1437, n_20818, n_20819);
  nand g40363 (n_15749, \data_stack_mem[1] [0], n_12808);
  or g40364 (n_15446, wc529, n_3673);
  not gc529 (wc529, n_14590);
  or g40365 (n_19039, n_1439, n_13900);
  or g40366 (n_15944, wc530, n_13788);
  not gc530 (wc530, \data_stack_mem[3] [1]);
  or g40367 (n_16001, wc531, n_13138);
  not gc531 (wc531, sh_reg_in[0]);
  or g40368 (n_15943, \data_stack_mem[3] [1], wc532);
  not gc532 (wc532, n_13788);
  nand g40369 (n_19044, n_14468, n_1439);
  or g40370 (n_16996, wc533, n_13770);
  not gc533 (wc533, \out_fifo[0][0] [1]);
  nand g40371 (n_16575, n_16569, n_16570);
  or g40372 (n_15372, wc534, n_15371);
  not gc534 (wc534, n_14151);
  nand g40373 (n_16573, n_16565, n_16566);
  or g40374 (n_17000, wc535, n_13405);
  not gc535 (wc535, \out_fifo[4][0] [1]);
  or g40375 (n_16568, wc536, n_13405);
  not gc536 (wc536, \out_fifo[4][2] [0]);
  or g40376 (n_16564, wc537, n_13770);
  not gc537 (wc537, \out_fifo[0][2] [0]);
  nand g40377 (n_17005, n_16997, n_16998);
  nand g40378 (n_17007, n_17001, n_17002);
  or g40379 (n_15135, n_15134, wc538);
  not gc538 (wc538, n_13764);
  or g40380 (n_16007, wc539, n_13138);
  not gc539 (wc539, sh_reg_in[1]);
  or g40381 (n_13107, wc540, n_15645);
  not gc540 (wc540, n_13816);
  nand g40382 (n_15840, \data_stack_mem[8] [6], n_12801);
  or g40383 (n_16013, wc541, n_13138);
  not gc541 (wc541, sh_reg_in[2]);
  nand g40384 (n_15834, \data_stack_mem[8] [0], n_12801);
  nand g40385 (n_19350, n_14546, n_14174);
  or g40386 (n_16019, wc542, n_13138);
  not gc542 (wc542, sh_reg_in[3]);
  or g40387 (n_17044, wc543, n_13770);
  not gc543 (wc543, \out_fifo[0][1] [0]);
  or g40388 (n_15743, wc544, n_13140);
  not gc544 (wc544, sh_reg_in[6]);
  or g40389 (n_16025, wc545, n_13138);
  not gc545 (wc545, sh_reg_in[4]);
  or g40390 (n_17048, wc546, n_13405);
  not gc546 (wc546, \out_fifo[4][1] [0]);
  or g40391 (n_14464, n_3673, wc547);
  not gc547 (wc547, n_15039);
  nand g40392 (n_20820, n_13400, n_1411);
  or g40393 (n_20821, n_13400, n_1411);
  nand g40394 (n_1427, n_20820, n_20821);
  nand g40395 (n_15828, \data_stack_mem[8] [1], n_12801);
  nand g40396 (n_16527, n_16521, n_16522);
  nand g40397 (n_15822, \data_stack_mem[8] [2], n_12801);
  nand g40398 (n_16525, n_16517, n_16518);
  or g40399 (n_15473, wc548, n_14194);
  not gc548 (wc548, n_14546);
  or g40400 (n_16520, wc549, n_13405);
  not gc549 (wc549, \out_fifo[4][1] [1]);
  or g40401 (n_16516, wc550, n_13770);
  not gc550 (wc550, \out_fifo[0][1] [1]);
  nand g40402 (n_15816, \data_stack_mem[8] [3], n_12801);
  or g40403 (n_15472, n_13989, n_14546);
  or g40404 (n_14465, n_12739, n_15075);
  or g40405 (n_15737, wc551, n_13140);
  not gc551 (wc551, sh_reg_in[5]);
  or g40406 (n_15990, wc552, n_13788);
  not gc552 (wc552, n_37);
  nand g40407 (n_16479, n_16473, n_16474);
  or g40408 (n_15731, wc553, n_13140);
  not gc553 (wc553, sh_reg_in[3]);
  nand g40409 (n_16477, n_16469, n_16470);
  nand g40410 (n_17053, n_17045, n_17046);
  or g40411 (n_16472, wc554, n_13405);
  not gc554 (wc554, \out_fifo[4][1] [2]);
  or g40412 (n_16468, wc555, n_13770);
  not gc555 (wc555, \out_fifo[0][1] [2]);
  nand g40413 (n_15276, n_15274, n_15275);
  or g40414 (n_15725, wc556, n_13140);
  not gc556 (wc556, sh_reg_in[0]);
  or g40415 (n_15719, wc557, n_13140);
  not gc557 (wc557, sh_reg_in[7]);
  nand g40416 (n_15620, n_14467, n_4344);
  nand g40417 (n_16431, n_16425, n_16426);
  or g40418 (n_16283, \data_stack_mem[2] [2], wc558);
  not gc558 (wc558, n_12683);
  or g40419 (n_16031, wc559, n_13138);
  not gc559 (wc559, sh_reg_in[5]);
  nand g40420 (n_17055, n_17049, n_17050);
  or g40421 (n_16037, wc560, n_13138);
  not gc560 (wc560, sh_reg_in[6]);
  or g40422 (n_18552, n_18550, wc561);
  not gc561 (wc561, \data_stack_mem[8] [4]);
  or g40423 (n_17092, wc562, n_13770);
  not gc562 (wc562, \out_fifo[0][1] [8]);
  or g40424 (n_17096, wc563, n_13405);
  not gc563 (wc563, \out_fifo[4][1] [8]);
  nand g40425 (n_17101, n_17093, n_17094);
  or g40426 (n_16043, wc564, n_13138);
  not gc564 (wc564, sh_reg_in[7]);
  nand g40427 (n_18555, n_14519, n_1433);
  nand g40428 (n_16429, n_16421, n_16422);
  nand g40429 (n_17103, n_17097, n_17098);
  or g40430 (n_16424, wc565, n_13405);
  not gc565 (wc565, \out_fifo[4][1] [3]);
  or g40431 (n_16420, wc566, n_13770);
  not gc566 (wc566, \out_fifo[0][1] [3]);
  or g40432 (n_17140, wc567, n_13770);
  not gc567 (wc567, \out_fifo[0][1] [7]);
  or g40433 (n_17144, wc568, n_13405);
  not gc568 (wc568, \out_fifo[4][1] [7]);
  nand g40434 (n_17149, n_17141, n_17142);
  nand g40435 (n_15810, \data_stack_mem[8] [5], n_12801);
  nand g40436 (n_16383, n_16377, n_16378);
  nand g40437 (n_17151, n_17145, n_17146);
  nand g40438 (n_15804, \data_stack_mem[8] [4], n_12801);
  nand g40439 (n_15798, \data_stack_mem[8] [7], n_12801);
  nand g40440 (n_16381, n_16373, n_16374);
  nand g40441 (n_5807, n_16049, n_16050);
  nand g40442 (n_15791, \data_stack_mem[1] [7], n_12808);
  or g40443 (n_16376, wc569, n_13405);
  not gc569 (wc569, \out_fifo[4][1] [4]);
  nand g40444 (n_5791, n_16055, n_16056);
  or g40445 (n_16372, wc570, n_13770);
  not gc570 (wc570, \out_fifo[0][1] [4]);
  or g40446 (n_17188, wc571, n_13770);
  not gc571 (wc571, \out_fifo[0][1] [6]);
  nand g40447 (n_5391, n_16061, n_16062);
  or g40448 (n_17192, wc572, n_13405);
  not gc572 (wc572, \out_fifo[4][1] [6]);
  or g40449 (n_14517, n_3673, wc573);
  not gc573 (wc573, n_15093);
  nand g40450 (n_17197, n_17189, n_17190);
  nand g40451 (n_17199, n_17193, n_17194);
  nand g40452 (n_16335, n_16329, n_16330);
  or g40453 (n_13106, n_14086, wc574);
  not gc574 (wc574, n_13608);
  nand g40454 (n_16333, n_16325, n_16326);
  or g40455 (n_13110, wc575, n_14086);
  not gc575 (wc575, n_14131);
  or g40456 (n_16328, wc576, n_13405);
  not gc576 (wc576, \out_fifo[4][1] [5]);
  or g40457 (n_16324, wc577, n_13770);
  not gc577 (wc577, \out_fifo[0][1] [5]);
  nand g40458 (n_5603, n_16277, n_16278);
  nand g40459 (n_5315, n_16271, n_16272);
  or g40460 (n_17236, wc578, n_13405);
  not gc578 (wc578, \out_fifo[4][0] [4]);
  or g40461 (n_14518, n_12739, n_14874);
  or g40462 (n_17239, wc579, n_13770);
  not gc579 (wc579, \out_fifo[0][0] [4]);
  nand g40463 (n_17245, n_17237, n_17238);
  nand g40464 (n_16264, n_16259, n_16260);
  nand g40465 (n_17247, n_17241, n_17242);
  nand g40466 (n_16262, n_16255, n_16256);
  or g40467 (n_15950, n_13812, n_14153);
  or g40468 (n_16257, wc580, n_13405);
  not gc580 (wc580, \out_fifo[4][0] [0]);
  or g40469 (n_16253, wc581, n_13770);
  not gc581 (wc581, \out_fifo[0][0] [0]);
  or g40470 (n_17284, wc582, n_13405);
  not gc582 (wc582, \out_fifo[4][0] [5]);
  or g40471 (n_17287, wc583, n_13770);
  not gc583 (wc583, \out_fifo[0][0] [5]);
  nand g40472 (n_17293, n_17285, n_17286);
  nand g40473 (n_17295, n_17289, n_17290);
  nand g40474 (n_5319, n_17303, n_17304);
  nand g40475 (n_5607, n_17309, n_17310);
  nand g40476 (n_5535, n_16067, n_16068);
  nand g40477 (n_5099, n_17324, n_17325);
  nand g40478 (n_5387, n_17330, n_17331);
  or g40479 (n_18313, n_1429, n_13900);
  nand g40480 (n_5531, n_17336, n_17337);
  nand g40481 (n_5459, n_17342, n_17343);
  nand g40482 (n_5243, n_17348, n_17349);
  nand g40483 (n_5103, n_16073, n_16074);
  nand g40484 (n_5171, n_17354, n_17355);
  nand g40485 (n_18318, n_14539, n_1429);
  or g40486 (n_15713, wc584, n_13140);
  not gc584 (wc584, sh_reg_in[4]);
  or g40487 (n_15707, wc585, n_13140);
  not gc585 (wc585, sh_reg_in[2]);
  or g40488 (n_15951, wc586, n_13764);
  not gc586 (wc586, n_13812);
  nand g40489 (n_19368, n_14544, n_14172);
  or g40490 (n_13108, wc587, n_15624);
  not gc587 (wc587, n_14137);
  or g40491 (n_15464, n_14194, n_14544);
  or g40492 (n_15463, wc588, n_13989);
  not gc588 (wc588, n_14544);
  or g40493 (n_16175, wc589, n_13137);
  not gc589 (wc589, sh_reg_in[7]);
  or g40494 (n_15701, wc590, n_13140);
  not gc590 (wc590, sh_reg_in[1]);
  nand g40495 (n_15696, \data_stack_mem[7] [2], n_13105);
  or g40496 (n_16169, wc591, n_13137);
  not gc591 (wc591, sh_reg_in[6]);
  nand g40497 (n_5175, n_16079, n_16080);
  nand g40498 (n_15690, \data_stack_mem[7] [3], n_13105);
  or g40499 (n_16163, wc592, n_13137);
  not gc592 (wc592, sh_reg_in[5]);
  nand g40500 (n_5463, n_16085, n_16086);
  nand g40501 (n_16289, \data_stack_mem[2] [2], n_12606);
  nand g40502 (n_15684, \data_stack_mem[7] [0], n_13105);
  nand g40503 (n_5247, n_16091, n_16092);
  or g40504 (n_16157, wc593, n_13137);
  not gc593 (wc593, sh_reg_in[4]);
  or g40505 (n_14537, n_3673, wc594);
  not gc594 (wc594, n_15111);
  nand g40506 (n_15264, n_15262, n_15263);
  nand g40507 (n_15678, \data_stack_mem[7] [6], n_13105);
  or g40508 (n_16151, wc595, n_13137);
  not gc595 (wc595, sh_reg_in[3]);
  nand g40509 (n_4088, n_15965, n_15966);
  nand g40510 (n_5008, n_15536, n_15537);
  or g40511 (n_16145, wc596, n_13137);
  not gc596 (wc596, sh_reg_in[2]);
  nand g40512 (n_15672, \data_stack_mem[7] [1], n_13105);
  nand g40513 (n_15666, \data_stack_mem[7] [7], n_13105);
  or g40514 (n_16139, wc597, n_13137);
  not gc597 (wc597, sh_reg_in[1]);
  nand g40515 (n_5016, n_13139, n_15558);
  nand g40516 (n_15660, \data_stack_mem[7] [5], n_13105);
  or g40517 (n_14538, n_12739, n_14913);
  or g40518 (n_16133, wc598, n_13137);
  not gc598 (wc598, sh_reg_in[0]);
  nand g40519 (n_5795, n_16127, n_16128);
  nand g40520 (n_5803, n_16121, n_16122);
  nand g40521 (n_5779, n_16115, n_16116);
  or g40522 (n_13111, n_15630, wc599);
  not gc599 (wc599, n_13608);
  or g40523 (n_15021, n_15020, wc600);
  not gc600 (wc600, n_14237);
  or g40524 (n_17315, wc601, n_13812);
  not gc601 (wc601, \data_stack_mem[3] [1]);
  nand g40525 (n_5799, n_16103, n_16104);
  or g40526 (n_17856, wc602, n_13183);
  not gc602 (wc602, n_14575);
  nand g40527 (n_5783, n_16109, n_16110);
  nand g40528 (n_15654, \data_stack_mem[7] [4], n_13105);
  nand g40529 (n_17928, \out_fifo[6][0] [1], n_12758);
  nand g40530 (n_17934, \out_fifo[0][0] [1], n_12756);
  nand g40531 (n_16098, \out_fifo[2][2] [0], n_12757);
  nand g40532 (n_17940, \out_fifo[1][0] [1], n_12760);
  or g40533 (n_16103, n_13831, n_12769);
  nand g40534 (n_16104, \out_fifo[5][2] [0], n_12762);
  or g40535 (n_15371, wc603, n_15370);
  not gc603 (wc603, n_14153);
  or g40536 (n_16109, n_13831, n_12768);
  nand g40537 (n_16110, \out_fifo[1][2] [0], n_12760);
  or g40538 (n_16999, wc604, n_13404);
  not gc604 (wc604, \out_fifo[7][0] [1]);
  nand g40539 (n_17946, \out_fifo[5][0] [1], n_12762);
  or g40540 (n_17001, wc605, n_13406);
  not gc605 (wc605, \out_fifo[5][0] [1]);
  or g40541 (n_17002, wc606, n_13407);
  not gc606 (wc606, \out_fifo[6][0] [1]);
  or g40542 (n_13183, n_14808, n_12739);
  nand g40543 (n_17952, \out_fifo[2][0] [1], n_12757);
  nand g40544 (n_19113, \out_fifo[2][1] [2], n_12757);
  nand g40545 (n_19119, \out_fifo[2][1] [3], n_12757);
  nand g40546 (n_19125, \out_fifo[4][0] [8], n_12759);
  nand g40547 (n_19131, \out_fifo[6][0] [8], n_12758);
  nand g40548 (n_19137, \out_fifo[0][0] [8], n_12756);
  nand g40549 (n_19143, \out_fifo[1][0] [8], n_12760);
  nand g40550 (n_17958, \out_fifo[3][0] [1], n_12761);
  or g40551 (n_15134, n_15133, wc607);
  not gc607 (wc607, n_12917);
  or g40552 (n_15851, wc608, n_13135);
  not gc608 (wc608, sh_reg_in[1]);
  or g40553 (n_15845, wc609, n_13135);
  not gc609 (wc609, sh_reg_in[0]);
  nand g40554 (n_17964, \out_fifo[7][0] [1], n_12755);
  or g40555 (n_15839, wc610, n_12803);
  not gc610 (wc610, sh_reg_in[6]);
  nand g40556 (n_18135, \out_fifo[4][0] [2], n_12759);
  nand g40557 (n_14553, n_14150, n_15375);
  nand g40558 (n_18141, \out_fifo[6][0] [2], n_12758);
  or g40559 (n_17043, wc611, n_13744);
  not gc611 (wc611, \out_fifo[3][1] [0]);
  nand g40560 (n_18147, \out_fifo[0][0] [2], n_12756);
  or g40561 (n_17045, wc612, n_13769);
  not gc612 (wc612, \out_fifo[1][1] [0]);
  nand g40562 (n_19149, \out_fifo[5][0] [8], n_12762);
  nand g40563 (n_19155, \out_fifo[3][0] [8], n_12761);
  nand g40564 (n_19161, \out_fifo[2][0] [8], n_12757);
  or g40565 (n_15020, n_15019, wc613);
  not gc613 (wc613, n_14294);
  or g40566 (n_17046, wc614, n_13768);
  not gc614 (wc614, \out_fifo[2][1] [0]);
  or g40567 (n_17047, wc615, n_13404);
  not gc615 (wc615, \out_fifo[7][1] [0]);
  nand g40568 (n_19167, \out_fifo[7][0] [8], n_12755);
  or g40569 (n_17049, wc616, n_13406);
  not gc616 (wc616, \out_fifo[5][1] [0]);
  or g40570 (n_20822, wc617, n_12929);
  not gc617 (wc617, n_13922);
  or g40571 (n_20823, n_13922, wc618);
  not gc618 (wc618, n_12929);
  nand g40572 (n_1411, n_20822, n_20823);
  or g40573 (n_15833, wc619, n_12803);
  not gc619 (wc619, sh_reg_in[0]);
  or g40574 (n_15827, wc620, n_12803);
  not gc620 (wc620, sh_reg_in[1]);
  or g40575 (n_15821, wc621, n_12803);
  not gc621 (wc621, sh_reg_in[2]);
  nand g40576 (n_14546, n_13920, n_15285);
  nand g40577 (n_19173, \out_fifo[7][1] [4], n_12755);
  nand g40578 (n_19179, \out_fifo[2][1] [4], n_12757);
  nand g40579 (n_18153, \out_fifo[1][0] [2], n_12760);
  nand g40580 (n_18159, \out_fifo[5][0] [2], n_12762);
  nand g40581 (n_18165, \out_fifo[3][0] [2], n_12761);
  nand g40582 (n_18171, \out_fifo[2][0] [2], n_12757);
  or g40583 (n_17050, wc622, n_13407);
  not gc622 (wc622, \out_fifo[6][1] [0]);
  nand g40584 (n_18177, \out_fifo[7][0] [2], n_12755);
  or g40585 (n_16115, n_13831, n_12767);
  nand g40586 (n_16116, \out_fifo[0][2] [0], n_12756);
  nand g40587 (n_15989, n_14237, n_1345);
  or g40588 (n_16121, n_13831, n_12766);
  nand g40589 (n_16122, \out_fifo[6][2] [0], n_12758);
  nand g40590 (n_18327, \out_fifo[4][0] [3], n_12759);
  or g40591 (n_16127, n_13831, n_12765);
  nand g40592 (n_16128, \out_fifo[4][2] [0], n_12759);
  nand g40593 (n_18333, \out_fifo[6][0] [3], n_12758);
  nand g40594 (n_18339, \out_fifo[0][0] [3], n_12756);
  or g40595 (n_14913, wc623, n_14912);
  not gc623 (wc623, n_14130);
  nand g40596 (n_18345, \out_fifo[1][0] [3], n_12760);
  or g40597 (n_15274, n_15273, wc624);
  not gc624 (wc624, n_3793);
  nand g40598 (n_18351, \out_fifo[5][0] [3], n_12762);
  nand g40599 (n_18357, \out_fifo[3][0] [3], n_12761);
  nand g40600 (n_18363, \out_fifo[2][0] [3], n_12757);
  nand g40601 (n_18369, \out_fifo[7][0] [3], n_12755);
  nand g40602 (n_18438, \out_fifo[4][0] [4], n_12759);
  nand g40603 (n_18444, \out_fifo[6][0] [4], n_12758);
  nand g40604 (n_18450, \out_fifo[0][0] [4], n_12756);
  nand g40605 (n_18456, \out_fifo[1][0] [4], n_12760);
  or g40606 (n_15111, n_15110, wc625);
  not gc625 (wc625, n_13767);
  or g40607 (n_16097, n_13831, n_12774);
  nand g40608 (n_16092, \out_fifo[2][2] [8], n_12757);
  or g40609 (n_16091, n_12774, status[7]);
  nand g40610 (n_16086, \out_fifo[5][2] [8], n_12762);
  or g40611 (n_16085, n_12769, status[7]);
  nand g40612 (n_16080, \out_fifo[1][2] [8], n_12760);
  nand g40613 (n_18462, \out_fifo[5][0] [4], n_12762);
  nand g40614 (n_18468, \out_fifo[3][0] [4], n_12761);
  nand g40615 (n_18474, \out_fifo[2][0] [4], n_12757);
  nand g40616 (n_14539, n_14150, n_15342);
  nand g40617 (n_18480, \out_fifo[7][0] [4], n_12755);
  or g40618 (n_16181, wc626, n_13832);
  not gc626 (wc626, sh_reg_in[7]);
  nand g40619 (n_19185, \out_fifo[3][1] [4], n_12761);
  nand g40620 (n_18564, \out_fifo[4][0] [5], n_12759);
  or g40621 (n_16187, wc627, n_13832);
  not gc627 (wc627, sh_reg_in[6]);
  nand g40622 (n_18570, \out_fifo[6][0] [5], n_12758);
  nand g40623 (n_18576, \out_fifo[0][0] [5], n_12756);
  or g40624 (n_16193, wc628, n_13832);
  not gc628 (wc628, sh_reg_in[3]);
  nand g40625 (n_19311, \out_fifo[0][1] [0], n_12756);
  nand g40626 (n_20824, n_13402, n_1413);
  or g40627 (n_20825, n_13402, n_1413);
  nand g40628 (n_1429, n_20824, n_20825);
  or g40629 (n_16199, wc629, n_13832);
  not gc629 (wc629, sh_reg_in[2]);
  or g40630 (n_16079, n_12768, status[7]);
  nand g40631 (n_18582, \out_fifo[1][0] [5], n_12760);
  or g40632 (n_16205, wc630, n_13832);
  not gc630 (wc630, sh_reg_in[1]);
  nand g40633 (n_16074, \out_fifo[0][2] [8], n_12756);
  or g40634 (n_15653, wc631, n_13139);
  not gc631 (wc631, sh_reg_in[4]);
  or g40635 (n_16211, wc632, n_13832);
  not gc632 (wc632, sh_reg_in[0]);
  or g40636 (n_16073, n_12767, status[7]);
  nand g40637 (n_16068, \out_fifo[6][2] [8], n_12758);
  or g40638 (n_16217, wc633, n_13832);
  not gc633 (wc633, sh_reg_in[5]);
  nand g40639 (n_5012, n_15299, n_15300);
  nand g40640 (n_19317, \out_fifo[1][1] [0], n_12760);
  or g40641 (n_16223, wc634, n_13832);
  not gc634 (wc634, sh_reg_in[4]);
  nand g40642 (n_19323, \out_fifo[5][1] [0], n_12762);
  nand g40643 (n_19329, \out_fifo[3][1] [0], n_12761);
  nand g40644 (n_19335, \out_fifo[2][1] [0], n_12757);
  or g40645 (n_13770, out_fifo_read_pointer[0], n_15993);
  nand g40646 (n_19341, \out_fifo[7][1] [0], n_12755);
  or g40647 (n_16254, wc635, n_13769);
  not gc635 (wc635, \out_fifo[1][0] [0]);
  or g40648 (n_16255, wc636, n_13768);
  not gc636 (wc636, \out_fifo[2][0] [0]);
  or g40649 (n_16256, wc637, n_13404);
  not gc637 (wc637, \out_fifo[7][0] [0]);
  or g40650 (n_15750, wc638, n_12806);
  not gc638 (wc638, sh_reg_in[0]);
  or g40651 (n_13405, out_fifo_read_pointer[0], n_15996);
  or g40652 (n_15263, n_15261, wc639);
  not gc639 (wc639, n_3793);
  or g40653 (n_15756, wc640, n_12806);
  not gc640 (wc640, sh_reg_in[1]);
  or g40654 (n_16258, wc641, n_13406);
  not gc641 (wc641, \out_fifo[5][0] [0]);
  or g40655 (n_16259, wc642, n_13407);
  not gc642 (wc642, \out_fifo[6][0] [0]);
  or g40656 (n_16260, wc643, n_13744);
  not gc643 (wc643, \out_fifo[3][0] [0]);
  or g40657 (n_15624, wc644, n_13967);
  not gc644 (wc644, n_14132);
  or g40658 (n_15659, wc645, n_13139);
  not gc645 (wc645, sh_reg_in[5]);
  or g40659 (n_15630, wc646, n_13452);
  not gc646 (wc646, n_15629);
  or g40660 (n_15815, wc647, n_12803);
  not gc647 (wc647, sh_reg_in[3]);
  or g40661 (n_15665, wc648, n_13139);
  not gc648 (wc648, sh_reg_in[7]);
  nand g40662 (n_18588, \out_fifo[5][0] [5], n_12762);
  or g40663 (n_14874, wc649, n_14873);
  not gc649 (wc649, n_14145);
  nand g40664 (n_16271, \out_fifo[3][2] [1], n_12761);
  or g40665 (n_16272, n_139, n_13244);
  nand g40666 (n_18594, \out_fifo[3][0] [5], n_12761);
  nand g40667 (n_16277, \out_fifo[7][2] [1], n_12755);
  or g40668 (n_16278, n_139, n_13242);
  nand g40669 (n_18600, \out_fifo[2][0] [5], n_12757);
  or g40670 (n_16323, wc650, n_13744);
  not gc650 (wc650, \out_fifo[3][1] [5]);
  nand g40671 (n_18606, \out_fifo[7][0] [5], n_12755);
  or g40672 (n_16325, wc651, n_13769);
  not gc651 (wc651, \out_fifo[1][1] [5]);
  or g40673 (n_16326, wc652, n_13768);
  not gc652 (wc652, \out_fifo[2][1] [5]);
  or g40674 (n_16327, wc653, n_13404);
  not gc653 (wc653, \out_fifo[7][1] [5]);
  nand g40675 (n_18681, \out_fifo[4][0] [6], n_12759);
  or g40676 (n_16329, wc654, n_13406);
  not gc654 (wc654, \out_fifo[5][1] [5]);
  or g40677 (n_16330, wc655, n_13407);
  not gc655 (wc655, \out_fifo[6][1] [5]);
  nand g40678 (n_15621, n_15618, n_15619);
  nand g40679 (n_18687, \out_fifo[6][0] [6], n_12758);
  nand g40680 (n_18693, \out_fifo[0][0] [6], n_12756);
  nand g40681 (n_18699, \out_fifo[1][0] [6], n_12760);
  nand g40682 (n_18705, \out_fifo[5][0] [6], n_12762);
  or g40683 (n_14467, n_15318, wc656);
  not gc656 (wc656, n_3902);
  nand g40684 (n_18711, \out_fifo[3][0] [6], n_12761);
  or g40685 (n_15093, n_15092, wc657);
  not gc657 (wc657, n_13766);
  or g40686 (n_16067, n_12766, status[7]);
  or g40687 (n_16371, wc658, n_13744);
  not gc658 (wc658, \out_fifo[3][1] [4]);
  nand g40688 (n_16062, \out_fifo[4][2] [8], n_12759);
  nand g40689 (n_18717, \out_fifo[2][0] [6], n_12757);
  or g40690 (n_16374, wc659, n_13768);
  not gc659 (wc659, \out_fifo[2][1] [4]);
  or g40691 (n_16375, wc660, n_13404);
  not gc660 (wc660, \out_fifo[7][1] [4]);
  or g40692 (n_16061, n_12765, status[7]);
  or g40693 (n_16377, wc661, n_13406);
  not gc661 (wc661, \out_fifo[5][1] [4]);
  or g40694 (n_16378, wc662, n_13407);
  not gc662 (wc662, \out_fifo[6][1] [4]);
  nand g40695 (n_18723, \out_fifo[7][0] [6], n_12755);
  nand g40696 (n_16056, \out_fifo[3][2] [0], n_12761);
  or g40697 (n_16055, n_13831, n_12772);
  nand g40698 (n_16050, \out_fifo[7][2] [0], n_12755);
  or g40699 (n_16049, n_13831, n_12775);
  nand g40700 (n_18792, \out_fifo[4][0] [7], n_12759);
  nand g40701 (n_14519, n_14150, n_15336);
  nand g40702 (n_18798, \out_fifo[6][0] [7], n_12758);
  nand g40703 (n_18804, \out_fifo[0][0] [7], n_12756);
  or g40704 (n_16419, wc663, n_13744);
  not gc663 (wc663, \out_fifo[3][1] [3]);
  nand g40705 (n_18810, \out_fifo[1][0] [7], n_12760);
  or g40706 (n_16421, wc664, n_13769);
  not gc664 (wc664, \out_fifo[1][1] [3]);
  or g40707 (n_16422, wc665, n_13768);
  not gc665 (wc665, \out_fifo[2][1] [3]);
  or g40708 (n_16423, wc666, n_13404);
  not gc666 (wc666, \out_fifo[7][1] [3]);
  nand g40709 (n_18816, \out_fifo[5][0] [7], n_12762);
  or g40710 (n_16425, wc667, n_13406);
  not gc667 (wc667, \out_fifo[5][1] [3]);
  or g40711 (n_16426, wc668, n_13407);
  not gc668 (wc668, \out_fifo[6][1] [3]);
  nand g40712 (n_18822, \out_fifo[3][0] [7], n_12761);
  nand g40713 (n_18828, \out_fifo[2][0] [7], n_12757);
  or g40714 (n_15762, wc669, n_12806);
  not gc669 (wc669, sh_reg_in[2]);
  or g40715 (n_12801, n_13939, wc670);
  not gc670 (wc670, n_15633);
  or g40716 (n_18550, n_1433, n_13900);
  nand g40717 (n_18834, \out_fifo[7][0] [7], n_12755);
  nand g40718 (n_18873, \out_fifo[4][1] [1], n_12759);
  nand g40719 (n_18879, \out_fifo[6][1] [1], n_12758);
  nand g40720 (n_12683, n_15605, n_15606);
  or g40721 (n_16467, wc671, n_13744);
  not gc671 (wc671, \out_fifo[3][1] [2]);
  nand g40722 (n_18885, \out_fifo[0][1] [1], n_12756);
  or g40723 (n_16469, wc672, n_13769);
  not gc672 (wc672, \out_fifo[1][1] [2]);
  or g40724 (n_16470, wc673, n_13768);
  not gc673 (wc673, \out_fifo[2][1] [2]);
  or g40725 (n_16471, wc674, n_13404);
  not gc674 (wc674, \out_fifo[7][1] [2]);
  nand g40726 (n_18891, \out_fifo[1][1] [1], n_12760);
  or g40727 (n_16473, wc675, n_13406);
  not gc675 (wc675, \out_fifo[5][1] [2]);
  or g40728 (n_16474, wc676, n_13407);
  not gc676 (wc676, \out_fifo[6][1] [2]);
  nand g40729 (n_18897, \out_fifo[5][1] [1], n_12762);
  nand g40730 (n_18903, \out_fifo[2][1] [1], n_12757);
  nand g40731 (n_18906, \out_fifo[6][1] [7], n_12758);
  or g40732 (n_15671, wc677, n_13139);
  not gc677 (wc677, sh_reg_in[1]);
  or g40733 (n_15965, wc678, n_4056);
  not gc678 (wc678, n_14477);
  or g40734 (n_15966, n_14477, wc679);
  not gc679 (wc679, n_4056);
  or g40735 (n_15677, wc680, n_13139);
  not gc680 (wc680, sh_reg_in[6]);
  or g40736 (n_15075, wc681, n_15074);
  not gc681 (wc681, n_14127);
  or g40737 (n_15683, wc682, n_13139);
  not gc682 (wc682, sh_reg_in[0]);
  or g40738 (n_15645, wc683, n_13967);
  not gc683 (wc683, n_15644);
  or g40739 (n_16515, wc684, n_13744);
  not gc684 (wc684, \out_fifo[3][1] [1]);
  or g40740 (n_15689, wc685, n_13139);
  not gc685 (wc685, sh_reg_in[3]);
  nand g40741 (n_12606, n_15527, n_19371);
  nand g40742 (n_15536, n_14569, rst_n);
  or g40743 (n_15768, wc686, n_12806);
  not gc686 (wc686, sh_reg_in[3]);
  or g40744 (n_16517, wc687, n_13769);
  not gc687 (wc687, \out_fifo[1][1] [1]);
  or g40745 (n_16518, wc688, n_13768);
  not gc688 (wc688, \out_fifo[2][1] [1]);
  or g40746 (n_16519, wc689, n_13404);
  not gc689 (wc689, \out_fifo[7][1] [1]);
  or g40747 (n_15774, wc690, n_12806);
  not gc690 (wc690, sh_reg_in[4]);
  or g40748 (n_16521, wc691, n_13406);
  not gc691 (wc691, \out_fifo[5][1] [1]);
  or g40749 (n_16522, wc692, n_13407);
  not gc692 (wc692, \out_fifo[6][1] [1]);
  nand g40750 (n_19191, \out_fifo[5][1] [4], n_12762);
  or g40751 (n_12808, n_13939, wc693);
  not gc693 (wc693, n_13816);
  nand g40752 (n_19197, \out_fifo[1][1] [4], n_12760);
  nand g40753 (n_19203, \out_fifo[0][1] [4], n_12756);
  nand g40754 (n_18909, \out_fifo[6][1] [8], n_12758);
  or g40755 (n_17091, wc694, n_13744);
  not gc694 (wc694, \out_fifo[3][1] [8]);
  nand g40756 (n_18912, \out_fifo[6][1] [6], n_12758);
  or g40757 (n_15039, n_15038, wc695);
  not gc695 (wc695, n_13765);
  or g40758 (n_17093, wc696, n_13769);
  not gc696 (wc696, \out_fifo[1][1] [8]);
  or g40759 (n_16563, wc697, n_13744);
  not gc697 (wc697, \out_fifo[3][2] [0]);
  nand g40760 (n_14468, n_14150, n_15321);
  or g40761 (n_16565, wc698, n_13769);
  not gc698 (wc698, \out_fifo[1][2] [0]);
  or g40762 (n_16566, wc699, n_13768);
  not gc699 (wc699, \out_fifo[2][2] [0]);
  or g40763 (n_16567, wc700, n_13404);
  not gc700 (wc700, \out_fifo[7][2] [0]);
  or g40764 (n_17094, wc701, n_13768);
  not gc701 (wc701, \out_fifo[2][1] [8]);
  or g40765 (n_16569, wc702, n_13406);
  not gc702 (wc702, \out_fifo[5][2] [0]);
  or g40766 (n_16570, wc703, n_13407);
  not gc703 (wc703, \out_fifo[6][2] [0]);
  or g40767 (n_17095, wc704, n_13404);
  not gc704 (wc704, \out_fifo[7][1] [8]);
  nand g40768 (n_18915, \out_fifo[6][1] [5], n_12758);
  or g40769 (n_17097, wc705, n_13406);
  not gc705 (wc705, \out_fifo[5][1] [8]);
  or g40770 (n_17098, wc706, n_13407);
  not gc706 (wc706, \out_fifo[6][1] [8]);
  nand g40771 (n_18918, \out_fifo[7][1] [8], n_12755);
  nand g40772 (n_19209, \out_fifo[6][1] [4], n_12758);
  nand g40773 (n_20826, n_13401, n_1423);
  or g40774 (n_20827, n_13401, n_1423);
  nand g40775 (n_1439, n_20826, n_20827);
  or g40776 (n_15780, wc707, n_12806);
  not gc707 (wc707, sh_reg_in[5]);
  nand g40777 (n_19215, \out_fifo[4][1] [4], n_12759);
  or g40778 (n_16611, wc708, n_13744);
  not gc708 (wc708, \out_fifo[3][2] [8]);
  nand g40779 (n_18921, \out_fifo[7][1] [5], n_12755);
  or g40780 (n_16613, wc709, n_13769);
  not gc709 (wc709, \out_fifo[1][2] [8]);
  or g40781 (n_16614, wc710, n_13768);
  not gc710 (wc710, \out_fifo[2][2] [8]);
  or g40782 (n_16615, wc711, n_13404);
  not gc711 (wc711, \out_fifo[7][2] [8]);
  nand g40783 (n_18924, \out_fifo[7][1] [6], n_12755);
  or g40784 (n_16617, wc712, n_13406);
  not gc712 (wc712, \out_fifo[5][2] [8]);
  or g40785 (n_16618, wc713, n_13407);
  not gc713 (wc713, \out_fifo[6][2] [8]);
  nand g40786 (n_18927, \out_fifo[7][1] [7], n_12755);
  nand g40787 (n_18930, \out_fifo[5][1] [5], n_12762);
  nand g40788 (n_18933, \out_fifo[5][1] [8], n_12762);
  or g40789 (n_17139, wc714, n_13744);
  not gc714 (wc714, \out_fifo[3][1] [7]);
  nand g40790 (n_18936, \out_fifo[5][1] [7], n_12762);
  or g40791 (n_17141, wc715, n_13769);
  not gc715 (wc715, \out_fifo[1][1] [7]);
  or g40792 (n_17142, wc716, n_13768);
  not gc716 (wc716, \out_fifo[2][1] [7]);
  or g40793 (n_17143, wc717, n_13404);
  not gc717 (wc717, \out_fifo[7][1] [7]);
  nand g40794 (n_18939, \out_fifo[5][1] [6], n_12762);
  or g40795 (n_16659, wc718, n_13744);
  not gc718 (wc718, \out_fifo[3][2] [1]);
  or g40796 (n_17145, wc719, n_13406);
  not gc719 (wc719, \out_fifo[5][1] [7]);
  or g40797 (n_16661, wc720, n_13769);
  not gc720 (wc720, \out_fifo[1][2] [1]);
  or g40798 (n_16662, wc721, n_13768);
  not gc721 (wc721, \out_fifo[2][2] [1]);
  or g40799 (n_16663, wc722, n_13404);
  not gc722 (wc722, \out_fifo[7][2] [1]);
  or g40800 (n_17146, wc723, n_13407);
  not gc723 (wc723, \out_fifo[6][1] [7]);
  or g40801 (n_16665, wc724, n_13406);
  not gc724 (wc724, \out_fifo[5][2] [1]);
  or g40802 (n_16666, wc725, n_13407);
  not gc725 (wc725, \out_fifo[6][2] [1]);
  nand g40803 (n_18942, \out_fifo[4][1] [8], n_12759);
  nand g40804 (n_18945, \out_fifo[4][1] [6], n_12759);
  nand g40805 (n_18948, \out_fifo[4][1] [7], n_12759);
  nand g40806 (n_18951, \out_fifo[4][1] [5], n_12759);
  nand g40807 (n_20828, n_13977, n_1403);
  or g40808 (n_20829, n_13977, n_1403);
  nand g40809 (n_1419, n_20828, n_20829);
  nand g40810 (n_18954, \out_fifo[0][1] [8], n_12756);
  or g40811 (n_15809, wc726, n_12803);
  not gc726 (wc726, sh_reg_in[5]);
  nand g40812 (n_14512, n_14150, n_15333);
  or g40813 (n_15803, wc727, n_12803);
  not gc727 (wc727, sh_reg_in[4]);
  or g40814 (n_16707, wc728, n_13744);
  not gc728 (wc728, \out_fifo[3][2] [9]);
  or g40815 (n_15797, wc729, n_12803);
  not gc729 (wc729, sh_reg_in[7]);
  or g40816 (n_15935, wc730, n_13134);
  not gc730 (wc730, sh_reg_in[4]);
  or g40817 (n_16709, wc731, n_13769);
  not gc731 (wc731, \out_fifo[1][2] [9]);
  or g40818 (n_16710, wc732, n_13768);
  not gc732 (wc732, \out_fifo[2][2] [9]);
  or g40819 (n_16711, wc733, n_13404);
  not gc733 (wc733, \out_fifo[7][2] [9]);
  or g40820 (n_15792, wc734, n_12806);
  not gc734 (wc734, sh_reg_in[7]);
  or g40821 (n_16713, wc735, n_13406);
  not gc735 (wc735, \out_fifo[5][2] [9]);
  or g40822 (n_16714, wc736, n_13407);
  not gc736 (wc736, \out_fifo[6][2] [9]);
  nand g40823 (n_18957, \out_fifo[0][1] [6], n_12756);
  or g40824 (n_17187, wc737, n_13744);
  not gc737 (wc737, \out_fifo[3][1] [6]);
  nand g40825 (n_18960, \out_fifo[0][1] [7], n_12756);
  or g40826 (n_17189, wc738, n_13769);
  not gc738 (wc738, \out_fifo[1][1] [6]);
  nand g40827 (n_18963, \out_fifo[0][1] [5], n_12756);
  or g40828 (n_17190, wc739, n_13768);
  not gc739 (wc739, \out_fifo[2][1] [6]);
  or g40829 (n_17191, wc740, n_13404);
  not gc740 (wc740, \out_fifo[7][1] [6]);
  nand g40830 (n_18966, \out_fifo[1][1] [7], n_12760);
  nand g40831 (n_18969, \out_fifo[1][1] [5], n_12760);
  or g40832 (n_16755, wc741, n_13744);
  not gc741 (wc741, \out_fifo[3][0] [8]);
  or g40833 (n_17193, wc742, n_13406);
  not gc742 (wc742, \out_fifo[5][1] [6]);
  or g40834 (n_16757, wc743, n_13769);
  not gc743 (wc743, \out_fifo[1][0] [8]);
  or g40835 (n_16758, wc744, n_13768);
  not gc744 (wc744, \out_fifo[2][0] [8]);
  or g40836 (n_17194, wc745, n_13407);
  not gc745 (wc745, \out_fifo[6][1] [6]);
  or g40837 (n_16759, wc746, n_13404);
  not gc746 (wc746, \out_fifo[7][0] [8]);
  nand g40838 (n_18972, \out_fifo[1][1] [8], n_12760);
  nand g40839 (n_18975, \out_fifo[1][1] [6], n_12760);
  or g40840 (n_14586, n_15429, n_12739);
  nand g40841 (n_18978, \out_fifo[3][1] [8], n_12761);
  nand g40842 (n_18981, \out_fifo[3][1] [5], n_12761);
  nand g40843 (n_18984, \out_fifo[3][1] [6], n_12761);
  nand g40844 (n_18987, \out_fifo[3][1] [7], n_12761);
  or g40845 (n_16761, wc747, n_13406);
  not gc747 (wc747, \out_fifo[5][0] [8]);
  or g40846 (n_16762, wc748, n_13407);
  not gc748 (wc748, \out_fifo[6][0] [8]);
  nand g40847 (n_18990, \out_fifo[2][1] [7], n_12757);
  or g40848 (n_14086, wc749, n_13452);
  not gc749 (wc749, n_15594);
  or g40849 (n_15434, wc750, n_3673);
  not gc750 (wc750, n_14587);
  nand g40850 (n_18993, \out_fifo[2][1] [6], n_12757);
  or g40851 (n_15435, n_14125, wc751);
  not gc751 (wc751, n_14172);
  or g40852 (n_15929, wc752, n_13134);
  not gc752 (wc752, sh_reg_in[5]);
  or g40853 (n_15923, wc753, n_13134);
  not gc753 (wc753, sh_reg_in[7]);
  or g40854 (n_15917, wc754, n_13134);
  not gc754 (wc754, sh_reg_in[6]);
  or g40855 (n_13137, n_14131, n_37);
  or g40856 (n_16803, wc755, n_13744);
  not gc755 (wc755, \out_fifo[3][0] [7]);
  or g40857 (n_17235, wc756, n_13407);
  not gc756 (wc756, \out_fifo[6][0] [4]);
  or g40858 (n_16805, wc757, n_13769);
  not gc757 (wc757, \out_fifo[1][0] [7]);
  or g40859 (n_16806, wc758, n_13768);
  not gc758 (wc758, \out_fifo[2][0] [7]);
  or g40860 (n_16807, wc759, n_13404);
  not gc759 (wc759, \out_fifo[7][0] [7]);
  nand g40861 (n_18996, \out_fifo[2][1] [8], n_12757);
  or g40862 (n_16809, wc760, n_13406);
  not gc760 (wc760, \out_fifo[5][0] [7]);
  or g40863 (n_16810, wc761, n_13407);
  not gc761 (wc761, \out_fifo[6][0] [7]);
  or g40864 (n_13138, n_14131, n_13942);
  or g40865 (n_17237, wc762, n_13404);
  not gc762 (wc762, \out_fifo[7][0] [4]);
  or g40866 (n_17238, wc763, n_13406);
  not gc763 (wc763, \out_fifo[5][0] [4]);
  nand g40867 (n_19221, \out_fifo[3][1] [2], n_12761);
  or g40868 (n_17240, wc764, n_13769);
  not gc764 (wc764, \out_fifo[1][0] [4]);
  or g40869 (n_17241, wc765, n_13768);
  not gc765 (wc765, \out_fifo[2][0] [4]);
  or g40870 (n_17242, wc766, n_13744);
  not gc766 (wc766, \out_fifo[3][0] [4]);
  nand g40871 (n_19227, \out_fifo[7][1] [2], n_12755);
  nand g40872 (n_20830, n_13952, n_1399);
  or g40873 (n_20831, n_13952, n_1399);
  nand g40874 (n_1415, n_20830, n_20831);
  or g40875 (n_16851, wc767, n_13744);
  not gc767 (wc767, \out_fifo[3][0] [6]);
  nand g40876 (n_19233, \out_fifo[3][1] [3], n_12761);
  or g40877 (n_16853, wc768, n_13769);
  not gc768 (wc768, \out_fifo[1][0] [6]);
  or g40878 (n_16854, wc769, n_13768);
  not gc769 (wc769, \out_fifo[2][0] [6]);
  or g40879 (n_16855, wc770, n_13404);
  not gc770 (wc770, \out_fifo[7][0] [6]);
  nand g40880 (n_14532, n_14150, n_15339);
  or g40881 (n_16857, wc771, n_13406);
  not gc771 (wc771, \out_fifo[5][0] [6]);
  or g40882 (n_16858, wc772, n_13407);
  not gc772 (wc772, \out_fifo[6][0] [6]);
  nand g40883 (n_19239, \out_fifo[7][1] [3], n_12755);
  nand g40884 (n_19251, \out_fifo[4][0] [0], n_12759);
  nand g40885 (n_19257, \out_fifo[6][0] [0], n_12758);
  nand g40886 (n_19263, \out_fifo[0][0] [0], n_12756);
  or g40887 (n_14588, n_15159, wc773);
  not gc773 (wc773, n_13803);
  or g40888 (n_15441, n_14125, wc774);
  not gc774 (wc774, n_14171);
  nand g40889 (n_19269, \out_fifo[1][0] [0], n_12760);
  nand g40890 (n_19275, \out_fifo[5][0] [0], n_12762);
  nand g40891 (n_14544, n_13918, n_15282);
  nand g40892 (n_19281, \out_fifo[3][0] [0], n_12761);
  nand g40893 (n_19287, \out_fifo[2][0] [0], n_12757);
  nand g40894 (n_5615, n_15542, n_15543);
  or g40895 (n_15695, wc775, n_13139);
  not gc775 (wc775, sh_reg_in[2]);
  or g40896 (n_15786, wc776, n_12806);
  not gc776 (wc776, sh_reg_in[6]);
  or g40897 (n_15558, n_15556, wc777);
  not gc777 (wc777, rst_n);
  or g40898 (n_17283, wc778, n_13407);
  not gc778 (wc778, \out_fifo[6][0] [5]);
  or g40899 (n_17453, n_14126, n_4054);
  or g40900 (n_17285, wc779, n_13404);
  not gc779 (wc779, \out_fifo[7][0] [5]);
  or g40901 (n_17286, wc780, n_13406);
  not gc780 (wc780, \out_fifo[5][0] [5]);
  or g40902 (n_16899, wc781, n_13744);
  not gc781 (wc781, \out_fifo[3][0] [3]);
  or g40903 (n_14589, n_12739, n_15198);
  or g40904 (n_16901, wc782, n_13769);
  not gc782 (wc782, \out_fifo[1][0] [3]);
  or g40905 (n_16902, wc783, n_13768);
  not gc783 (wc783, \out_fifo[2][0] [3]);
  or g40906 (n_16903, wc784, n_13404);
  not gc784 (wc784, \out_fifo[7][0] [3]);
  or g40907 (n_15911, wc785, n_13134);
  not gc785 (wc785, sh_reg_in[1]);
  or g40908 (n_16905, wc786, n_13406);
  not gc786 (wc786, \out_fifo[5][0] [3]);
  or g40909 (n_16906, wc787, n_13407);
  not gc787 (wc787, \out_fifo[6][0] [3]);
  or g40910 (n_13140, data_stack_pointer[3], n_15495);
  or g40911 (n_15905, wc788, n_13134);
  not gc788 (wc788, sh_reg_in[0]);
  or g40912 (n_15899, wc789, n_13134);
  not gc789 (wc789, sh_reg_in[2]);
  or g40913 (n_13109, n_13939, n_15639);
  or g40914 (n_15893, wc790, n_13134);
  not gc790 (wc790, sh_reg_in[3]);
  or g40915 (n_17288, wc791, n_13769);
  not gc791 (wc791, \out_fifo[1][0] [5]);
  or g40916 (n_15887, wc792, n_13135);
  not gc792 (wc792, sh_reg_in[7]);
  or g40917 (n_17289, wc793, n_13768);
  not gc793 (wc793, \out_fifo[2][0] [5]);
  or g40918 (n_17290, wc794, n_13744);
  not gc794 (wc794, \out_fifo[3][0] [5]);
  or g40919 (n_16947, wc795, n_13744);
  not gc795 (wc795, \out_fifo[3][0] [2]);
  or g40920 (n_13105, n_13452, wc796);
  not gc796 (wc796, n_15648);
  or g40921 (n_16949, wc797, n_13769);
  not gc797 (wc797, \out_fifo[1][0] [2]);
  or g40922 (n_16950, wc798, n_13768);
  not gc798 (wc798, \out_fifo[2][0] [2]);
  or g40923 (n_16951, wc799, n_13404);
  not gc799 (wc799, \out_fifo[7][0] [2]);
  or g40924 (n_16373, wc800, n_13769);
  not gc800 (wc800, \out_fifo[1][1] [4]);
  or g40925 (n_16953, wc801, n_13406);
  not gc801 (wc801, \out_fifo[5][0] [2]);
  or g40926 (n_16954, wc802, n_13407);
  not gc802 (wc802, \out_fifo[6][0] [2]);
  nand g40927 (n_19293, \out_fifo[7][0] [0], n_12755);
  nand g40928 (n_18999, \out_fifo[2][1] [5], n_12757);
  nand g40929 (n_19005, \out_fifo[3][1] [1], n_12761);
  nand g40930 (n_19011, \out_fifo[7][1] [1], n_12755);
  nand g40931 (n_19053, \out_fifo[4][1] [2], n_12759);
  nand g40932 (n_19059, \out_fifo[4][1] [3], n_12759);
  nand g40933 (n_19299, \out_fifo[4][1] [0], n_12759);
  or g40934 (n_17303, n_12772, status[7]);
  nand g40935 (n_20832, n_13969, n_1405);
  or g40936 (n_20833, n_13969, n_1405);
  nand g40937 (n_1421, n_20832, n_20833);
  nand g40938 (n_17304, \out_fifo[3][2] [8], n_12761);
  nand g40939 (n_14495, n_14150, n_15330);
  nand g40940 (n_19305, \out_fifo[6][1] [0], n_12758);
  or g40941 (n_17309, n_12775, status[7]);
  nand g40942 (n_17310, \out_fifo[7][2] [8], n_12755);
  nand g40943 (n_19065, \out_fifo[6][1] [2], n_12758);
  nand g40944 (n_19071, \out_fifo[6][1] [3], n_12758);
  nand g40945 (n_5619, n_12772, n_17319);
  nand g40946 (n_17324, n_12756, \out_fifo[0][2] [1]);
  or g40947 (n_17325, n_12921, n_13244);
  nand g40948 (n_19077, \out_fifo[0][1] [2], n_12756);
  nand g40949 (n_17330, n_12759, \out_fifo[4][2] [1]);
  or g40950 (n_17331, n_12921, n_13242);
  nand g40951 (n_19083, \out_fifo[0][1] [3], n_12756);
  nand g40952 (n_17336, n_12758, \out_fifo[6][2] [1]);
  or g40953 (n_17337, n_12854, n_13242);
  or g40954 (n_14591, n_15252, n_12739);
  nand g40955 (n_19089, \out_fifo[1][1] [2], n_12760);
  nand g40956 (n_17342, n_12762, \out_fifo[5][2] [1]);
  or g40957 (n_17343, n_12847, n_13242);
  nand g40958 (n_19095, \out_fifo[1][1] [3], n_12760);
  or g40959 (n_14590, n_15210, wc803);
  not gc803 (wc803, n_13970);
  or g40960 (n_15447, n_14125, wc804);
  not gc804 (wc804, n_13774);
  or g40961 (n_15881, wc805, n_13135);
  not gc805 (wc805, sh_reg_in[6]);
  or g40962 (n_15875, wc806, n_13135);
  not gc806 (wc806, sh_reg_in[5]);
  or g40963 (n_15869, wc807, n_13135);
  not gc807 (wc807, sh_reg_in[4]);
  or g40964 (n_15863, wc808, n_13135);
  not gc808 (wc808, sh_reg_in[3]);
  or g40965 (n_15857, wc809, n_13135);
  not gc809 (wc809, sh_reg_in[2]);
  nand g40966 (n_17348, n_12757, \out_fifo[2][2] [1]);
  or g40967 (n_17349, n_12854, n_13244);
  nand g40968 (n_19101, \out_fifo[5][1] [2], n_12762);
  nand g40969 (n_17354, n_12760, \out_fifo[1][2] [1]);
  or g40970 (n_16995, wc810, n_13744);
  not gc810 (wc810, \out_fifo[3][0] [1]);
  or g40971 (n_17355, n_12847, n_13244);
  or g40972 (n_16997, wc811, n_13769);
  not gc811 (wc811, \out_fifo[1][0] [1]);
  or g40973 (n_16998, wc812, n_13768);
  not gc812 (wc812, \out_fifo[2][0] [1]);
  nand g40974 (n_19107, \out_fifo[5][1] [3], n_12762);
  nand g40975 (n_17922, \out_fifo[4][0] [1], n_12759);
  or g40976 (n_15495, data_stack_pointer[0], n_15494);
  or g40977 (n_13996, n_15000, wc813);
  not gc813 (wc813, n_11331);
  nand g40978 (n_19371, n_14232, n_4056);
  or g40979 (n_15648, wc814, n_13449);
  not gc814 (wc814, n_14556);
  or g40980 (n_15629, wc815, n_13449);
  not gc815 (wc815, n_13942);
  or g40981 (n_13139, data_stack_pointer[3], n_15555);
  or g40982 (n_14574, n_14916, wc816);
  not gc816 (wc816, n_3634);
  nand g40983 (n_15556, n_14571, data_stack_pointer[3]);
  nand g40984 (n_15542, n_14570, rst_n);
  or g40985 (n_12739, sh_reg_in[1], n_14766);
  nand g40986 (n_5611, n_15515, n_15516);
  or g40987 (n_4054, wc817, n_14997);
  not gc817 (wc817, n_14140);
  or g40988 (n_12803, n_15498, wc818);
  not gc818 (wc818, data_stack_pointer[3]);
  or g40989 (n_14808, n_14807, wc819);
  not gc819 (wc819, \data_stack_mem[0] [0]);
  nand g40990 (n_13967, n_15452, n_15453);
  nand g40991 (n_14569, n_15386, n_15387);
  or g40992 (n_15262, n_14142, n_11312);
  or g40993 (n_15261, n_13428, wc820);
  not gc820 (wc820, n_11312);
  or g40994 (n_15300, data_stack_pointer[2], n_13608);
  nand g40995 (n_15282, n_13794, n_11312);
  nand g40996 (n_14477, n_15326, n_15327);
  nand g40997 (n_5031, n_14732, n_14733);
  or g40998 (n_5027, wc821, n_14700);
  not gc821 (wc821, n_14699);
  nand g40999 (n_17319, n_14557, out_fifo_write_pointer[2]);
  or g41000 (n_13244, out_fifo_write_pointer[2], n_14167);
  or g41001 (n_12772, n_857, wc822);
  not gc822 (wc822, rst_n);
  or g41002 (n_12775, n_817, wc823);
  not gc823 (wc823, rst_n);
  or g41003 (n_13242, n_14167, wc824);
  not gc824 (wc824, out_fifo_write_pointer[2]);
  nand g41004 (n_12761, n_13995, n_13940);
  nand g41005 (n_12755, n_13982, n_13940);
  or g41006 (n_13407, n_12753, n_12734);
  or g41007 (n_15019, n_15018, wc825);
  not gc825 (wc825, n_14246);
  or g41008 (n_13404, n_12732, n_12753);
  or g41009 (n_13406, n_12753, n_12733);
  or g41010 (n_14131, data_stack_pointer[0], n_13449);
  or g41011 (n_15594, wc826, n_13449);
  not gc826 (wc826, n_37);
  or g41012 (n_12767, n_13961, wc827);
  not gc827 (wc827, rst_n);
  or g41013 (n_12769, n_13956, wc828);
  not gc828 (wc828, rst_n);
  or g41014 (n_12774, n_13951, wc829);
  not gc829 (wc829, rst_n);
  or g41015 (n_12768, n_13949, wc830);
  not gc830 (wc830, rst_n);
  or g41016 (n_12766, n_13947, wc831);
  not gc831 (wc831, rst_n);
  or g41017 (n_12765, n_13946, wc832);
  not gc832 (wc832, rst_n);
  nand g41018 (n_13939, n_15453, n_13808);
  or g41019 (n_15605, \data_stack_mem[2] [1], wc833);
  not gc833 (wc833, n_14266);
  or g41020 (n_13832, n_37, n_13608);
  nand g41021 (n_15318, n_15316, n_15317);
  or g41022 (n_14912, wc834, n_14911);
  not gc834 (wc834, n_14152);
  or g41023 (n_15618, n_15617, wc835);
  not gc835 (wc835, n_13784);
  or g41024 (n_15619, n_13825, n_14266);
  or g41025 (n_13744, n_12732, n_12754);
  or g41026 (n_13769, n_12754, n_12733);
  or g41027 (n_13768, n_12754, n_12734);
  or g41028 (n_4342, wc836, n_14970);
  not gc836 (wc836, n_14140);
  or g41029 (n_12806, data_stack_pointer[2], n_15501);
  or g41030 (n_15273, n_13428, n_119);
  or g41031 (n_15275, n_14142, wc837);
  not gc837 (wc837, n_119);
  or g41032 (n_15110, n_15109, wc838);
  not gc838 (wc838, n_13402);
  nand g41033 (n_1345, n_15479, n_15480);
  or g41034 (n_14150, wc839, n_12777);
  not gc839 (wc839, n_11331);
  or g41035 (n_15342, \data_stack_mem[8] [2], n_12777);
  nand g41036 (n_15285, n_13795, n_119);
  or g41037 (n_20834, wc840, n_12896);
  not gc840 (wc840, n_1379);
  or g41038 (n_20835, n_1379, wc841);
  not gc841 (wc841, n_12896);
  nand g41039 (n_13922, n_20834, n_20835);
  or g41040 (n_15375, \data_stack_mem[8] [1], n_12777);
  or g41041 (n_13135, n_13903, n_15494);
  or g41042 (n_15133, n_15132, wc842);
  not gc842 (wc842, n_13400);
  or g41043 (n_20836, wc843, n_12871);
  not gc843 (wc843, n_13901);
  or g41044 (n_20837, n_13901, wc844);
  not gc844 (wc844, n_12871);
  nand g41045 (n_1413, n_20836, n_20837);
  or g41046 (n_13450, n_11331, n_15000);
  or g41047 (n_13900, n_12777, n_11331);
  or g41048 (n_15370, n_15368, n_15369);
  or g41049 (n_15210, n_15209, wc845);
  not gc845 (wc845, n_13950);
  or g41050 (n_15330, \data_stack_mem[8] [6], n_12777);
  nand g41051 (n_20838, n_13971, n_1389);
  or g41052 (n_20839, n_13971, n_1389);
  nand g41053 (n_1405, n_20838, n_20839);
  or g41054 (n_15993, out_fifo_read_pointer[1], n_12754);
  or g41055 (n_13134, data_stack_pointer[3], n_15498);
  or g41056 (n_15996, out_fifo_read_pointer[1], n_12753);
  or g41057 (n_15198, wc846, n_15197);
  not gc846 (wc846, n_14126);
  or g41058 (n_15159, n_15158, wc847);
  not gc847 (wc847, n_13980);
  or g41059 (n_15339, \data_stack_mem[8] [3], n_12777);
  nand g41060 (n_20840, n_13975, n_1383);
  or g41061 (n_20841, n_13975, n_1383);
  nand g41062 (n_1399, n_20840, n_20841);
  or g41063 (n_14125, wc848, n_3673);
  not gc848 (wc848, n_3793);
  or g41064 (n_14587, n_15147, wc849);
  not gc849 (wc849, n_13912);
  or g41065 (n_15429, n_15427, n_15428);
  or g41066 (n_14873, wc850, n_14872);
  not gc850 (wc850, n_14133);
  nand g41067 (n_12756, n_13995, n_15954);
  or g41068 (n_15333, \data_stack_mem[8] [5], n_12777);
  nand g41069 (n_12759, n_15954, n_13982);
  nand g41070 (n_20842, n_13976, n_1387);
  or g41071 (n_20843, n_13976, n_1387);
  nand g41072 (n_1403, n_20842, n_20843);
  nand g41073 (n_12758, n_13982, n_15957);
  nand g41074 (n_12757, n_15957, n_13995);
  nand g41075 (n_12762, n_13982, n_15960);
  nand g41076 (n_12760, n_15960, n_13995);
  or g41077 (n_20844, wc851, n_12861);
  not gc851 (wc851, n_13902);
  or g41078 (n_20845, n_13902, wc852);
  not gc852 (wc852, n_12861);
  nand g41079 (n_1423, n_20844, n_20845);
  or g41080 (n_15321, \data_stack_mem[8] [7], n_12777);
  or g41081 (n_15092, n_15091, wc853);
  not gc853 (wc853, n_13403);
  or g41082 (n_15038, n_15037, wc854);
  not gc854 (wc854, n_13401);
  or g41083 (n_15074, wc855, n_15073);
  not gc855 (wc855, n_14136);
  or g41084 (n_15336, \data_stack_mem[8] [4], n_12777);
  nand g41085 (n_20846, n_13403, n_1417);
  or g41086 (n_20847, n_13403, n_1417);
  nand g41087 (n_1433, n_20846, n_20847);
  or g41088 (n_15617, n_4344, n_12917);
  nand g41089 (n_13831, n_4634, status[7]);
  nand g41090 (n_14997, n_14995, n_14996);
  or g41091 (n_15317, wc856, n_13784);
  not gc856 (wc856, \data_stack_mem[2] [1]);
  nand g41092 (n_20848, n_13905, n_1385);
  or g41093 (n_20849, n_13905, n_1385);
  nand g41094 (n_1417, n_20848, n_20849);
  or g41095 (n_15316, \data_stack_mem[2] [1], wc857);
  not gc857 (wc857, n_13784);
  or g41096 (n_13449, n_15489, wc858);
  not gc858 (wc858, data_stack_pointer[1]);
  or g41097 (n_4343, wc859, n_14949);
  not gc859 (wc859, n_13986);
  or g41098 (n_15132, n_15131, wc860);
  not gc860 (wc860, n_12941);
  or g41099 (n_15000, n_3634, wc861);
  not gc861 (wc861, n_4634);
  or g41100 (n_20850, wc862, n_12862);
  not gc862 (wc862, n_1381);
  or g41101 (n_20851, n_1381, wc863);
  not gc863 (wc863, n_12862);
  nand g41102 (n_13901, n_20850, n_20851);
  nand g41103 (n_20852, n_13964, n_1367);
  or g41104 (n_20853, n_13964, n_1367);
  nand g41105 (n_1383, n_20852, n_20853);
  nand g41106 (n_5643, n_12738, n_15567);
  or g41107 (n_15326, n_13811, n_13825);
  nand g41108 (n_5651, n_12738, n_15522);
  or g41109 (n_12753, wc864, n_12738);
  not gc864 (wc864, out_fifo_read_pointer[2]);
  nand g41110 (n_14557, n_14147, n_13940);
  or g41111 (n_15073, n_15071, n_15072);
  or g41112 (n_15158, n_15157, wc865);
  not gc865 (wc865, n_13975);
  or g41113 (n_20854, wc866, n_12941);
  not gc866 (wc866, n_13904);
  or g41114 (n_20855, n_13904, wc867);
  not gc867 (wc867, n_12941);
  nand g41115 (n_1379, n_20854, n_20855);
  or g41116 (n_14766, n_14765, wc868);
  not gc868 (wc868, sh_reg_in[0]);
  or g41117 (n_13608, sh_reg_in[8], n_15486);
  or g41118 (n_14911, n_14909, n_14910);
  or g41119 (n_15501, n_14137, n_1483);
  nand g41120 (n_15606, n_13784, n_4344);
  or g41121 (n_15543, wc869, n_14147);
  not gc869 (wc869, out_fifo_write_pointer[1]);
  or g41122 (n_15386, n_15384, wc870);
  not gc870 (wc870, data_stack_pointer[0]);
  or g41123 (n_15527, wc871, n_13811);
  not gc871 (wc871, \data_stack_mem[2] [1]);
  or g41124 (n_14733, n_14731, wc872);
  not gc872 (wc872, rst_n);
  or g41125 (n_15037, n_15036, wc873);
  not gc873 (wc873, n_14173);
  or g41126 (n_15197, n_15195, n_15196);
  or g41127 (n_12777, n_14143, wc874);
  not gc874 (wc874, n_4634);
  or g41128 (n_15109, n_15108, wc875);
  not gc875 (wc875, n_12869);
  nand g41129 (n_119, n_14667, n_19347);
  nand g41130 (n_5019, n_12738, n_15504);
  or g41131 (n_14732, out_fifo_read_pointer[2], n_14730);
  or g41132 (n_15555, n_13789, n_15554);
  or g41133 (n_20856, wc876, n_12870);
  not gc876 (wc876, n_1391);
  or g41134 (n_20857, n_1391, wc877);
  not gc877 (wc877, n_12870);
  nand g41135 (n_13902, n_20856, n_20857);
  or g41136 (n_15091, n_15090, wc878);
  not gc878 (wc878, n_12932);
  or g41137 (n_15018, n_15017, wc879);
  not gc879 (wc879, n_14209);
  or g41138 (n_15327, n_12917, wc880);
  not gc880 (wc880, n_13811);
  or g41139 (n_12754, out_fifo_read_pointer[2], n_12738);
  or g41140 (n_15480, wc881, n_13784);
  not gc881 (wc881, n_3902);
  nand g41141 (n_14570, n_12854, n_15390);
  nand g41142 (n_14916, n_14143, n_3637);
  or g41143 (n_14135, wc882, n_13817);
  not gc882 (wc882, n_4634);
  nand g41144 (n_15453, n_1483, rst_n);
  nand g41145 (n_20858, n_13970, n_1373);
  or g41146 (n_20859, n_13970, n_1373);
  nand g41147 (n_1389, n_20858, n_20859);
  or g41148 (n_15299, n_13808, wc883);
  not gc883 (wc883, n_13917);
  nand g41149 (n_14700, n_14697, n_14698);
  or g41150 (n_14571, n_13917, wc884);
  not gc884 (wc884, n_15393);
  nand g41151 (n_5635, n_12738, n_15507);
  nand g41152 (n_14970, n_14968, n_14969);
  or g41153 (n_4055, wc885, n_14937);
  not gc885 (wc885, n_13986);
  nand g41154 (n_20860, n_13966, n_1371);
  or g41155 (n_20861, n_13966, n_1371);
  nand g41156 (n_1387, n_20860, n_20861);
  or g41157 (n_15515, n_15514, wc886);
  not gc886 (wc886, rst_n);
  or g41158 (n_15494, n_13808, n_1483);
  or g41159 (n_15498, n_14132, n_1483);
  nand g41160 (n_5023, n_14705, n_14706);
  or g41161 (n_857, n_139, n_13215);
  not g41162 (n_20862, n_857);
  or g41163 (n_15252, n_15250, n_15251);
  or g41164 (n_817, n_139, n_13214);
  not g41165 (n_20863, n_817);
  nand g41166 (n_5004, n_15305, n_15306);
  or g41167 (n_15427, wc887, n_15424);
  not gc887 (wc887, n_15423);
  or g41168 (n_15209, n_15208, wc888);
  not gc888 (wc888, n_13978);
  or g41169 (n_15516, wc889, n_14147);
  not gc889 (wc889, out_fifo_write_pointer[0]);
  or g41170 (n_14807, n_14805, n_14806);
  nand g41171 (n_5647, n_12738, n_15564);
  or g41172 (n_14167, n_4634, n_15456);
  nand g41173 (n_11312, n_14820, n_19365);
  or g41174 (n_3673, sh_reg_in[0], n_14143);
  nand g41175 (n_13982, rst_n, n_13214);
  or g41176 (n_15369, wc890, n_15367);
  not gc890 (wc890, n_15366);
  or g41177 (n_15147, n_15146, wc891);
  not gc891 (wc891, n_13966);
  nand g41178 (n_13995, rst_n, n_13215);
  or g41179 (n_14872, n_14870, n_14871);
  or g41180 (n_17291, wc892, n_11);
  not gc892 (wc892, sh_reg_out[4]);
  or g41181 (n_17051, wc893, n_11);
  not gc893 (wc893, sh_reg_out[9]);
  or g41182 (n_14910, n_14907, n_14908);
  or g41183 (n_15387, data_stack_pointer[0], n_15385);
  or g41184 (n_16427, wc894, n_11);
  not gc894 (wc894, sh_reg_out[12]);
  or g41185 (n_20864, wc895, n_1353);
  not gc895 (wc895, n_13533);
  or g41186 (n_20865, n_13533, wc896);
  not gc896 (wc896, n_1353);
  nand g41187 (n_1385, n_20864, n_20865);
  or g41188 (n_16955, wc897, n_11);
  not gc897 (wc897, sh_reg_out[1]);
  or g41189 (n_15456, n_13925, wc898);
  not gc898 (wc898, sh_reg_in[8]);
  or g41190 (n_15384, data_stack_pointer[1], n_14168);
  nand g41191 (n_14147, rst_n, n_131);
  or g41192 (n_15306, wc899, n_14166);
  not gc899 (wc899, data_stack_pointer[0]);
  or g41193 (n_15131, n_15130, wc900);
  not gc900 (wc900, n_12929);
  or g41194 (n_16475, wc901, n_11);
  not gc901 (wc901, sh_reg_out[11]);
  or g41195 (n_15017, n_15016, wc902);
  not gc902 (wc902, n_14196);
  or g41196 (n_17243, wc903, n_11);
  not gc903 (wc903, sh_reg_out[3]);
  nand g41197 (n_20866, n_13950, n_1357);
  or g41198 (n_20867, n_13950, n_1357);
  nand g41199 (n_1373, n_20866, n_20867);
  or g41200 (n_15072, n_15069, n_15070);
  or g41201 (n_15486, n_13789, n_13925);
  nand g41202 (n_14937, n_14935, n_14936);
  or g41203 (n_12764, n_11331, n_3637);
  or g41204 (n_5631, n_14166, wc904);
  not gc904 (wc904, n_15309);
  or g41205 (n_13917, n_158, wc905);
  not gc905 (wc905, n_15279);
  or g41208 (n_14968, n_13992, n_14530);
  or g41209 (n_14697, n_12733, n_14164);
  or g41210 (n_16523, wc906, n_11);
  not gc906 (wc906, sh_reg_out[10]);
  nand g41211 (n_13452, n_14166, n_15483);
  or g41212 (n_20869, wc907, n_1349);
  not gc907 (wc907, n_13536);
  or g41213 (n_20870, n_13536, wc908);
  not gc908 (wc908, n_1349);
  nand g41214 (n_1381, n_20869, n_20870);
  nand g41215 (n_14949, n_14947, n_14948);
  or g41216 (n_15036, n_15035, wc909);
  not gc909 (wc909, n_12920);
  or g41217 (n_16379, wc910, n_11);
  not gc910 (wc910, sh_reg_out[13]);
  or g41218 (n_15567, wc911, n_11);
  not gc911 (wc911, n_14582);
  or g41219 (n_15305, n_13816, n_14168);
  or g41220 (n_16571, wc912, n_11);
  not gc912 (wc912, sh_reg_out[19]);
  or g41221 (n_14698, wc913, n_14163);
  not gc913 (wc913, out_fifo_read_pointer[1]);
  or g41222 (n_15250, n_15246, n_15247);
  or g41223 (n_20871, wc914, n_1359);
  not gc914 (wc914, n_13538);
  or g41224 (n_20872, n_13538, wc915);
  not gc915 (wc915, n_1359);
  nand g41225 (n_1391, n_20871, n_20872);
  or g41226 (n_14705, out_fifo_read_pointer[0], n_14164);
  or g41227 (n_15090, n_15089, wc916);
  not gc916 (wc916, n_12933);
  or g41228 (n_15564, wc917, n_11);
  not gc917 (wc917, n_14581);
  or g41229 (n_14969, wc918, n_14193);
  not gc918 (wc918, n_14530);
  or g41230 (n_16619, wc919, n_11);
  not gc919 (wc919, sh_reg_out[27]);
  or g41231 (n_4056, wc920, n_14961);
  not gc920 (wc920, n_14159);
  or g41232 (n_15554, n_14168, n_13808);
  or g41233 (n_17195, wc921, n_11);
  not gc921 (wc921, sh_reg_out[15]);
  or g41234 (n_15537, wc922, n_14166);
  not gc922 (wc922, data_stack_pointer[1]);
  or g41235 (n_12738, wc923, n_14180);
  not gc923 (wc923, n_14566);
  or g41236 (n_15522, n_15521, n_11);
  or g41237 (n_15489, sh_reg_in[8], n_13925);
  or g41238 (n_14143, wc924, n_13953);
  not gc924 (wc924, sh_reg_in[1]);
  or g41239 (n_20873, wc925, n_13764);
  not gc925 (wc925, n_1347);
  or g41240 (n_20874, n_1347, wc926);
  not gc926 (wc926, n_13764);
  nand g41241 (n_13904, n_20873, n_20874);
  or g41242 (n_16667, wc927, n_11);
  not gc927 (wc927, sh_reg_out[20]);
  nand g41243 (n_20875, n_13979, n_1355);
  or g41244 (n_20876, n_13979, n_1355);
  nand g41245 (n_1371, n_20875, n_20876);
  or g41246 (n_16331, wc928, n_11);
  not gc928 (wc928, sh_reg_out[14]);
  or g41247 (n_17147, wc929, n_11);
  not gc929 (wc929, sh_reg_out[16]);
  nand g41248 (n_19365, n_14526, n_14171);
  or g41249 (n_14765, wc930, n_13953);
  not gc930 (wc930, n_14764);
  or g41250 (n_15514, n_131, out_fifo_write_pointer[0]);
  or g41253 (n_16715, wc931, n_11);
  not gc931 (wc931, sh_reg_out[28]);
  nand g41256 (n_5628, n_14834, n_14835);
  or g41257 (n_15424, n_1083, wc932);
  not gc932 (wc932, n_15418);
  or g41260 (n_15507, sh_reg_out_bit_counter[0], n_11);
  or g41261 (n_15251, n_15248, n_15249);
  nand g41264 (n_19347, n_14530, n_14175);
  or g41265 (n_15208, n_15207, wc933);
  not gc933 (wc933, n_13971);
  or g41266 (n_15428, n_15425, n_15426);
  or g41267 (n_15108, n_15107, wc934);
  not gc934 (wc934, n_12898);
  or g41268 (n_17099, wc935, n_11);
  not gc935 (wc935, sh_reg_out[17]);
  or g41271 (n_15146, n_15145, wc936);
  not gc936 (wc936, n_13979);
  or g41272 (n_16763, wc937, n_11);
  not gc937 (wc937, sh_reg_out[7]);
  or g41273 (n_14871, n_14868, n_14869);
  or g41274 (n_14706, wc938, n_14163);
  not gc938 (wc938, out_fifo_read_pointer[0]);
  or g41275 (n_15504, wc939, n_11);
  not gc939 (wc939, dout_valid);
  or g41276 (n_16811, wc940, n_11);
  not gc940 (wc940, sh_reg_out[6]);
  or g41277 (n_14995, wc941, n_13992);
  not gc941 (wc941, n_14526);
  or g41278 (n_14996, n_14193, n_14526);
  nand g41279 (n_14731, n_14584, out_fifo_read_pointer[2]);
  nand g41280 (status[7], n_14593, n_4634);
  nand g41281 (n_20882, n_13980, n_1351);
  or g41282 (n_20883, n_13980, n_1351);
  nand g41283 (n_1367, n_20882, n_20883);
  or g41286 (n_14806, n_14803, n_14804);
  or g41287 (n_16859, wc942, n_11);
  not gc942 (wc942, sh_reg_out[5]);
  or g41290 (n_15157, n_15156, wc943);
  not gc943 (wc943, n_13965);
  or g41293 (n_14730, n_12732, n_14164);
  nand g41294 (n_15479, n_14246, n_1329);
  nand g41295 (n_5625, n_14165, n_14919);
  or g41296 (n_15195, wc944, n_15192);
  not gc944 (wc944, n_15191);
  or g41297 (n_15367, n_1075, wc945);
  not gc945 (wc945, n_15363);
  or g41298 (n_15390, n_12847, n_131);
  or g41299 (n_3634, n_19344, wc946);
  not gc946 (wc946, sh_reg_in[4]);
  or g41300 (n_1483, data_stack_pointer[1], n_15288);
  or g41301 (n_15196, n_15193, n_15194);
  or g41302 (n_13817, wc947, n_3637);
  not gc947 (wc947, n_11331);
  or g41303 (n_16907, wc948, n_11);
  not gc948 (wc948, sh_reg_out[2]);
  or g41304 (n_17003, wc949, n_11);
  not gc949 (wc949, sh_reg_out[0]);
  or g41305 (n_4344, wc950, n_14988);
  not gc950 (wc950, n_14159);
  nand g41306 (n_14163, rst_n, n_100);
  nand g41307 (n_14907, n_14901, n_14902);
  nand g41308 (n_20887, n_12933, n_1337);
  or g41309 (n_20888, n_12933, n_1337);
  nand g41310 (n_1353, n_20887, n_20888);
  or g41311 (n_20889, wc951, n_12932);
  not gc951 (wc951, n_13766);
  or g41312 (n_20890, n_13766, wc952);
  not gc952 (wc952, n_12932);
  nand g41313 (n_13533, n_20889, n_20890);
  or g41314 (n_14164, n_100, wc953);
  not gc953 (wc953, rst_n);
  nand g41315 (n_15071, n_15067, n_15068);
  or g41316 (n_14936, n_14934, wc954);
  not gc954 (wc954, n_3793);
  nand g41317 (n_15069, n_12779, n_15064);
  nand g41318 (n_15070, n_15065, n_15066);
  nand g41319 (n_20891, n_12872, n_12863);
  or g41320 (n_20892, n_12872, n_12863);
  nand g41321 (n_13905, n_20891, n_20892);
  or g41322 (n_3637, n_14757, wc955);
  not gc955 (wc955, sh_reg_in[5]);
  nand g41323 (n_15016, n_14302, n_15015);
  or g41324 (n_15035, n_15034, wc956);
  not gc956 (wc956, n_12870);
  nand g41325 (n_15483, n_14559, rst_n);
  or g41326 (n_20893, wc957, n_12920);
  not gc957 (wc957, n_13765);
  or g41327 (n_20894, n_13765, wc958);
  not gc958 (wc958, n_12920);
  nand g41328 (n_13538, n_20893, n_20894);
  nand g41329 (n_20895, n_12866, n_1343);
  or g41330 (n_20896, n_12866, n_1343);
  nand g41331 (n_1359, n_20895, n_20896);
  nand g41332 (n_14909, n_14905, n_14906);
  or g41333 (n_15089, n_15088, wc959);
  not gc959 (wc959, n_12872);
  nand g41334 (n_14166, rst_n, n_158);
  or g41335 (n_20897, wc960, n_13797);
  not gc960 (wc960, n_13912);
  or g41336 (n_20898, n_13912, wc961);
  not gc961 (wc961, n_13797);
  nand g41337 (n_1355, n_20897, n_20898);
  or g41338 (n_13953, sh_reg_in[4], n_14664);
  nand g41339 (n_1083, n_14585, n_13821);
  nand g41340 (n_15425, n_15419, n_15420);
  nand g41341 (n_11, n_14178, rst_n);
  nand g41342 (n_15426, n_15421, n_15422);
  nand g41343 (n_14526, n_13919, n_14751);
  or g41344 (n_15145, n_15144, wc962);
  not gc962 (wc962, n_13977);
  or g41345 (n_20899, wc963, n_13803);
  not gc963 (wc963, n_13911);
  or g41346 (n_20900, n_13911, wc964);
  not gc964 (wc964, n_13803);
  nand g41347 (n_1351, n_20899, n_20900);
  nand g41348 (n_14869, n_14864, n_14865);
  nand g41349 (n_15156, n_13952, n_13964);
  nand g41350 (n_14908, n_14903, n_14904);
  or g41351 (n_19344, n_13933, n_14664);
  nand g41352 (n_1329, n_14975, n_14976);
  or g41353 (n_15393, data_stack_pointer[2], n_4615);
  nand g41354 (n_14988, n_14986, n_14987);
  nand g41355 (n_15194, n_15189, n_15190);
  nand g41356 (n_14868, n_14862, n_14863);
  nand g41357 (n_14804, n_14799, n_14800);
  or g41358 (n_15385, n_4615, wc965);
  not gc965 (wc965, data_stack_pointer[1]);
  or g41359 (n_15288, n_158, sh_reg_in[8]);
  or g41360 (n_20901, wc966, n_13804);
  not gc966 (wc966, n_13978);
  or g41361 (n_20902, n_13978, wc967);
  not gc967 (wc967, n_13804);
  nand g41362 (n_1357, n_20901, n_20902);
  or g41363 (n_14834, sh_bit_cnt[2], n_14165);
  nand g41364 (n_15246, n_12780, n_15239);
  or g41365 (n_14947, n_14946, wc968);
  not gc968 (wc968, n_3793);
  nand g41366 (n_15247, n_15240, n_15241);
  or g41367 (n_13925, n_158, wc969);
  not gc969 (wc969, rst_n);
  nand g41368 (n_15248, n_15242, n_15243);
  nand g41369 (n_14961, n_14959, n_14960);
  nand g41370 (n_15207, n_13959, n_13969);
  nand g41371 (n_14870, n_14866, n_14867);
  nand g41372 (n_14919, n_14580, rst_n);
  nand g41373 (n_15368, n_15364, n_15365);
  or g41374 (n_14593, n_14742, n_12864);
  or g41375 (n_15107, n_15106, wc970);
  not gc970 (wc970, n_12871);
  nand g41376 (n_1075, n_14592, n_13825);
  nand g41377 (n_15130, n_14550, n_12896);
  nand g41378 (n_14530, n_13907, n_14754);
  or g41379 (n_20903, wc971, n_12917);
  not gc971 (wc971, n_13913);
  or g41380 (n_20904, n_13913, wc972);
  not gc972 (wc972, n_12917);
  nand g41381 (n_1347, n_20903, n_20904);
  nand g41382 (n_20905, n_12898, n_1333);
  or g41383 (n_20906, n_12898, n_1333);
  nand g41384 (n_1349, n_20905, n_20906);
  or g41385 (n_14168, n_158, n_4615);
  nand g41386 (n_14803, n_14797, n_14798);
  or g41387 (n_20907, wc973, n_12869);
  not gc973 (wc973, n_13767);
  or g41388 (n_20908, n_13767, wc974);
  not gc974 (wc974, n_12869);
  nand g41389 (n_13536, n_20907, n_20908);
  or g41390 (n_15279, wc975, n_4615);
  not gc975 (wc975, n_13789);
  or g41391 (n_14180, n_14178, wc976);
  not gc976 (wc976, rst_n);
  nand g41392 (n_15192, n_12827, n_15186);
  nand g41393 (n_14975, \data_stack_mem[0] [0], n_14294);
  or g41394 (n_4615, sh_reg_in[8], wc977);
  not gc977 (wc977, n_14594);
  nand g41395 (n_14581, n_13121, n_14922);
  nand g41396 (n_1333, n_14148, n_13986);
  nand g41397 (n_13913, n_14128, n_14826);
  or g41398 (n_14866, \data_stack_mem[4] [4], n_20);
  nand g41399 (n_14754, n_13792, n_11358);
  or g41400 (n_12896, n_3910, wc978);
  not gc978 (wc978, \data_stack_mem[6] [1]);
  nand g41401 (n_15309, sh_bit_cnt[3], n_14281);
  nand g41402 (n_14867, n_13918, n_13981);
  or g41403 (n_15363, \data_stack_mem[8] [1], n_11331);
  or g41404 (n_12871, n_3910, wc979);
  not gc979 (wc979, \data_stack_mem[6] [2]);
  or g41405 (n_14960, n_14958, wc980);
  not gc980 (wc980, n_3793);
  or g41406 (n_14798, \data_stack_mem[6] [0], n_3910);
  or g41407 (n_14959, n_13916, n_14128);
  nand g41408 (n_14742, n_14740, n_14741);
  nand g41409 (n_14592, n_14682, n_14159);
  or g41410 (n_15366, \data_stack_mem[4] [1], n_20);
  nand g41411 (n_15106, n_14536, n_12862);
  or g41412 (n_14800, \data_stack_mem[4] [0], n_20);
  or g41413 (n_15364, \data_stack_mem[6] [1], n_3910);
  nand g41414 (n_15249, n_15244, n_15245);
  or g41415 (n_15242, \data_stack_mem[4] [6], n_20);
  or g41416 (n_14948, n_14148, wc981);
  not gc981 (wc981, n_11358);
  or g41417 (n_15241, \data_stack_mem[8] [6], n_11331);
  or g41418 (n_14946, n_170, n_11358);
  or g41419 (n_14835, n_14833, wc982);
  not gc982 (wc982, rst_n);
  or g41420 (n_15240, \data_stack_mem[6] [6], n_3910);
  nand g41421 (n_12780, n_13938, n_14134);
  or g41422 (n_14863, \data_stack_mem[8] [4], n_11331);
  nand g41423 (n_13804, n_14144, n_14823);
  or g41424 (n_13969, wc983, n_3910);
  not gc983 (wc983, \data_stack_mem[6] [6]);
  or g41425 (n_14987, n_14985, wc984);
  not gc984 (wc984, n_3793);
  or g41426 (n_14165, n_14745, wc985);
  not gc985 (wc985, rst_n);
  or g41427 (n_14986, n_14128, n_13814);
  or g41428 (n_15190, \data_stack_mem[8] [3], n_11331);
  or g41429 (n_15189, \data_stack_mem[4] [3], n_20);
  nand g41430 (n_15193, n_15187, n_15188);
  or g41431 (n_14664, n_12864, sh_reg_in[5]);
  or g41432 (n_14805, wc986, n_14802);
  not gc986 (wc986, n_14801);
  nand g41433 (n_12827, n_14140, n_14820);
  or g41434 (n_15191, \data_stack_mem[6] [3], n_3910);
  or g41435 (n_14864, \data_stack_mem[6] [4], n_3910);
  nand g41436 (n_13911, n_13992, n_14817);
  nand g41437 (n_14580, n_14717, n_14718);
  or g41438 (n_13952, wc987, n_3910);
  not gc987 (wc987, \data_stack_mem[6] [3]);
  nand g41439 (n_15144, n_13958, n_13976);
  nand g41440 (n_14751, n_13793, n_11305);
  or g41441 (n_15421, \data_stack_mem[8] [5], n_11331);
  or g41442 (n_15419, \data_stack_mem[6] [5], n_3910);
  nand g41443 (n_14585, n_14160, n_14925);
  or g41444 (n_15423, \data_stack_mem[4] [5], n_20);
  nand g41445 (n_15088, n_14516, n_12863);
  or g41446 (n_12872, n_3910, wc988);
  not gc988 (wc988, \data_stack_mem[6] [4]);
  nand g41447 (n_13797, n_13989, n_14814);
  nand g41448 (n_15521, sh_reg_out_bit_counter[4], n_13121);
  or g41449 (n_13977, wc989, n_3910);
  not gc989 (wc989, \data_stack_mem[6] [5]);
  or g41450 (n_14196, wc990, n_3910);
  not gc990 (wc990, \data_stack_mem[6] [0]);
  or g41451 (n_14559, sh_reg_in[8], n_14655);
  nand g41452 (n_1343, n_13987, n_13898);
  or g41453 (n_12870, n_3910, wc991);
  not gc991 (wc991, \data_stack_mem[6] [7]);
  nand g41454 (n_15034, n_12861, n_12866);
  nand g41455 (n_14906, n_13919, n_13986);
  or g41456 (n_14905, \data_stack_mem[4] [2], n_20);
  or g41457 (n_14757, n_14184, n_12864);
  or g41458 (n_15066, \data_stack_mem[8] [7], n_11331);
  or g41459 (n_15065, \data_stack_mem[4] [7], n_20);
  nand g41460 (n_12779, n_13987, n_14811);
  or g41461 (n_14902, \data_stack_mem[8] [2], n_11331);
  or g41462 (n_15068, \data_stack_mem[6] [7], n_3910);
  or g41463 (n_14903, \data_stack_mem[6] [2], n_3910);
  or g41464 (n_14934, n_170, wc992);
  not gc992 (wc992, n_11305);
  nand g41465 (n_1337, n_14142, n_13981);
  or g41466 (n_100, n_14637, wc993);
  not gc993 (wc993, sh_reg_out_bit_counter[0]);
  or g41467 (n_14935, n_14148, n_11305);
  or g41468 (n_14637, sh_reg_out_bit_counter[4], n_14636);
  or g41469 (n_14799, \data_stack_mem[5] [0], n_3908);
  or g41470 (n_15365, \data_stack_mem[5] [1], n_3908);
  nand g41471 (n_11331, data_stack_pointer[3], n_14685);
  or g41472 (n_15245, \data_stack_mem[2] [6], wc994);
  not gc994 (wc994, n_3902);
  or g41473 (n_14801, \data_stack_mem[1] [0], wc995);
  not gc995 (wc995, n_3793);
  nand g41474 (n_14142, n_3793, n_13428);
  or g41475 (n_14901, \data_stack_mem[2] [2], wc996);
  not gc996 (wc996, n_3902);
  or g41476 (n_13981, wc997, n_3793);
  not gc997 (wc997, \data_stack_mem[0] [4]);
  nand g41477 (n_20, n_37, n_14688);
  or g41478 (n_15243, \data_stack_mem[5] [6], n_3908);
  or g41479 (n_14862, \data_stack_mem[2] [4], wc998);
  not gc998 (wc998, n_3902);
  or g41480 (n_14823, \data_stack_mem[0] [6], n_3793);
  or g41481 (n_12861, n_3908, wc999);
  not gc999 (wc999, \data_stack_mem[5] [7]);
  or g41482 (n_5622, n_14649, wc1000);
  not gc1000 (wc1000, rst_n);
  or g41483 (n_13971, n_3908, wc1001);
  not gc1001 (wc1001, \data_stack_mem[5] [6]);
  or g41484 (n_14594, n_14661, wc1002);
  not gc1002 (wc1002, data_stack_pointer[3]);
  or g41485 (n_15188, \data_stack_mem[5] [3], n_3908);
  nand g41486 (n_15015, \data_stack_mem[0] [0], n_3793);
  nand g41487 (n_14655, n_13948, n_14654);
  or g41488 (n_15064, \data_stack_mem[5] [7], n_3908);
  nand g41489 (n_14173, n_3793, n_14748);
  or g41490 (n_19361, n_14811, wc1003);
  not gc1003 (wc1003, n_3793);
  nand g41491 (n_14802, n_14795, n_14796);
  or g41492 (n_14209, wc1004, n_3908);
  not gc1004 (wc1004, \data_stack_mem[5] [0]);
  or g41493 (n_14126, \data_stack_mem[2] [3], wc1005);
  not gc1005 (wc1005, n_3902);
  or g41494 (n_14192, wc1006, n_1327);
  not gc1006 (wc1006, n_3793);
  or g41495 (n_15067, \data_stack_mem[2] [7], wc1007);
  not gc1007 (wc1007, n_3902);
  or g41496 (n_14718, wc1008, n_13806);
  not gc1008 (wc1008, sh_bit_cnt[2]);
  or g41497 (n_14865, \data_stack_mem[5] [4], n_3908);
  nand g41498 (n_13898, n_3793, n_1327);
  nand g41499 (n_14193, n_3793, n_1323);
  or g41500 (n_13987, wc1009, n_3793);
  not gc1009 (wc1009, \data_stack_mem[0] [7]);
  nand g41501 (n_3910, n_37, n_14545);
  or g41502 (n_14817, \data_stack_mem[0] [3], n_3793);
  or g41503 (n_13992, wc1010, n_1323);
  not gc1010 (wc1010, n_3793);
  nand g41504 (n_14582, n_13934, n_14721);
  or g41505 (n_14904, \data_stack_mem[5] [2], n_3908);
  or g41506 (n_14144, wc1011, n_1326);
  not gc1011 (wc1011, n_3793);
  nand g41507 (n_11305, n_14681, n_14682);
  nand g41508 (n_15639, n_15638, n_14137);
  or g41509 (n_14797, \data_stack_mem[2] [0], wc1012);
  not gc1012 (wc1012, n_3902);
  or g41510 (n_13975, n_3908, wc1013);
  not gc1013 (wc1013, \data_stack_mem[5] [3]);
  or g41511 (n_14159, wc1014, n_3793);
  not gc1014 (wc1014, \data_stack_mem[0] [1]);
  or g41512 (n_14134, wc1015, n_3793);
  not gc1015 (wc1015, \data_stack_mem[0] [6]);
  or g41513 (n_14745, wc1016, n_13806);
  not gc1016 (wc1016, sh_bit_cnt[3]);
  or g41514 (n_12864, sh_reg_in[7], n_14643);
  nand g41515 (n_14985, n_168, n_13814);
  nand g41516 (n_14833, sh_bit_cnt[2], n_13806);
  or g41517 (n_13986, wc1017, n_3793);
  not gc1017 (wc1017, \data_stack_mem[0] [2]);
  nand g41518 (n_11358, n_14676, n_19356);
  nand g41519 (n_14194, n_3793, n_1325);
  or g41520 (n_13989, wc1018, n_1325);
  not gc1018 (wc1018, n_3793);
  or g41521 (n_14140, wc1019, n_3793);
  not gc1019 (wc1019, \data_stack_mem[0] [3]);
  or g41522 (n_14128, wc1020, n_168);
  not gc1020 (wc1020, n_3793);
  or g41523 (n_12862, n_3908, wc1021);
  not gc1021 (wc1021, \data_stack_mem[5] [2]);
  or g41524 (n_15420, \data_stack_mem[5] [5], n_3908);
  nand g41525 (n_14958, n_13916, n_168);
  nand g41526 (n_14740, sh_reg_in[5], n_14184);
  or g41527 (n_14160, wc1022, n_3793);
  not gc1022 (wc1022, \data_stack_mem[0] [5]);
  nand g41528 (n_14922, sh_reg_out_bit_counter[3], n_13934);
  nand g41529 (n_14148, n_3793, n_170);
  or g41530 (n_14976, wc1023, n_13814);
  not gc1023 (wc1023, n_3793);
  or g41531 (n_14621, n_14627, n_14628);
  or g41532 (n_12863, n_3908, wc1024);
  not gc1024 (wc1024, \data_stack_mem[5] [4]);
  or g41533 (n_14814, \data_stack_mem[0] [5], n_3793);
  or g41534 (n_13976, n_3908, wc1025);
  not gc1025 (wc1025, \data_stack_mem[5] [5]);
  or g41535 (n_14826, \data_stack_mem[0] [1], n_3793);
  or g41536 (n_12929, n_3908, wc1026);
  not gc1026 (wc1026, \data_stack_mem[5] [1]);
  or g41537 (n_14636, sh_reg_out_bit_counter[3], n_14635);
  nand g41538 (n_13764, \data_stack_mem[3] [1], n_37);
  or g41539 (n_14685, data_stack_pointer[0], n_13932);
  or g41540 (n_14153, wc1027, \data_stack_mem[3] [1]);
  not gc1027 (wc1027, n_37);
  or g41541 (n_14137, n_13903, wc1028);
  not gc1028 (wc1028, rst_n);
  nand g41542 (n_13940, n_139, rst_n);
  or g41543 (n_14796, \data_stack_mem[3] [0], wc1029);
  not gc1029 (wc1029, n_37);
  nand g41544 (n_14583, n_13815, n_14658);
  nand g41545 (n_14237, \data_stack_mem[3] [0], n_37);
  or g41546 (n_14132, data_stack_pointer[2], n_13816);
  or g41547 (n_14688, data_stack_pointer[0], n_13948);
  nand g41548 (n_14649, n_13778, n_14648);
  or g41549 (n_14661, wc1030, n_13932);
  not gc1030 (wc1030, data_stack_pointer[0]);
  or g41550 (n_3902, wc1031, n_37);
  not gc1031 (wc1031, n_13789);
  or g41551 (n_14699, n_12734, wc1032);
  not gc1032 (wc1032, rst_n);
  or g41552 (n_14136, wc1033, \data_stack_mem[3] [7]);
  not gc1033 (wc1033, n_37);
  nand g41553 (n_13765, \data_stack_mem[3] [7], n_37);
  or g41554 (n_14654, data_stack_pointer[1], wc1034);
  not gc1034 (wc1034, n_14558);
  nand g41555 (n_14717, sh_bit_cnt[1], n_13778);
  nand g41556 (n_1327, n_14170, n_14673);
  nand g41557 (n_14721, sh_reg_out_bit_counter[2], n_13815);
  or g41558 (n_3793, data_stack_pointer[1], n_37);
  or g41559 (n_14643, sh_reg_in[6], n_14642);
  nand g41560 (n_168, n_14296, n_14676);
  nand g41561 (n_1325, n_14174, n_14670);
  nand g41562 (n_14741, sh_reg_in[4], n_13933);
  or g41563 (n_14133, wc1035, \data_stack_mem[3] [4]);
  not gc1035 (wc1035, n_37);
  nand g41564 (n_14628, n_14625, n_14626);
  nand g41565 (n_14627, n_14623, n_14624);
  nand g41566 (n_13766, \data_stack_mem[3] [4], n_37);
  or g41567 (n_15244, \data_stack_mem[3] [6], wc1036);
  not gc1036 (wc1036, n_37);
  nand g41568 (n_13950, \data_stack_mem[3] [6], n_37);
  or g41569 (n_15452, wc1037, n_13808);
  not gc1037 (wc1037, data_stack_pointer[3]);
  or g41570 (n_15187, \data_stack_mem[3] [3], wc1038);
  not gc1038 (wc1038, n_37);
  nand g41571 (n_14764, data_stack_pointer[3], n_13932);
  nand g41572 (n_1323, n_14175, n_14667);
  nand g41573 (n_13980, \data_stack_mem[3] [3], n_37);
  or g41574 (n_15422, \data_stack_mem[3] [5], wc1039);
  not gc1039 (wc1039, n_37);
  nand g41575 (n_15954, n_12921, rst_n);
  nand g41576 (n_13979, \data_stack_mem[3] [5], n_37);
  nand g41577 (n_15957, n_12854, rst_n);
  nand g41578 (n_15960, n_12847, rst_n);
  nand g41579 (n_3908, n_37, n_13948);
  or g41580 (n_14130, wc1040, \data_stack_mem[3] [2]);
  not gc1040 (wc1040, n_37);
  or g41581 (n_15638, wc1041, n_13816);
  not gc1041 (wc1041, data_stack_pointer[3]);
  or g41582 (n_15644, n_37, wc1042);
  not gc1042 (wc1042, rst_n);
  nand g41583 (n_13767, \data_stack_mem[3] [2], n_37);
  or g41584 (n_14681, n_13916, wc1043);
  not gc1043 (wc1043, n_14297);
  nand g41585 (n_19356, n_13814, n_14296);
  nand g41586 (n_14682, \data_stack_mem[0] [1], \data_stack_mem[1] [1]);
  or g41587 (n_14667, wc1044, \data_stack_mem[1] [3]);
  not gc1044 (wc1044, \data_stack_mem[0] [3]);
  nand g41588 (n_14820, \data_stack_mem[0] [3], \data_stack_mem[1] [3]);
  or g41589 (n_14670, wc1045, \data_stack_mem[1] [5]);
  not gc1045 (wc1045, \data_stack_mem[0] [5]);
  or g41590 (n_14676, wc1046, \data_stack_mem[1] [1]);
  not gc1046 (wc1046, \data_stack_mem[0] [1]);
  nand g41591 (n_14925, \data_stack_mem[0] [5], \data_stack_mem[1] [5]);
  or g41592 (n_14673, \data_stack_mem[0] [7], wc1047);
  not gc1047 (wc1047, \data_stack_mem[1] [7]);
  nand g41593 (n_14811, \data_stack_mem[0] [7], \data_stack_mem[1] [7]);
  or g41594 (n_14748, \data_stack_mem[0] [7], \data_stack_mem[1] [7]);
  or g41595 (n_14127, \data_stack_mem[7] [7], wc1048);
  not gc1048 (wc1048, data_stack_pointer[3]);
  or g41596 (n_14145, \data_stack_mem[7] [4], wc1049);
  not gc1049 (wc1049, data_stack_pointer[3]);
  or g41597 (n_14152, \data_stack_mem[7] [2], wc1050);
  not gc1050 (wc1050, data_stack_pointer[3]);
  or g41598 (n_14151, \data_stack_mem[7] [1], wc1051);
  not gc1051 (wc1051, data_stack_pointer[3]);
  or g41599 (n_14642, sh_reg_in[2], sh_reg_in[3]);
  or g41600 (n_14795, \data_stack_mem[7] [0], wc1052);
  not gc1052 (wc1052, data_stack_pointer[3]);
  or g41601 (n_15418, \data_stack_mem[7] [5], wc1053);
  not gc1053 (wc1053, data_stack_pointer[3]);
  or g41602 (n_15186, \data_stack_mem[7] [3], wc1054);
  not gc1054 (wc1054, data_stack_pointer[3]);
  or g41603 (n_15239, \data_stack_mem[7] [6], wc1055);
  not gc1055 (wc1055, data_stack_pointer[3]);
  nand g41604 (n_139, out_fifo_write_pointer[0],
       out_fifo_write_pointer[1]);
  or g41605 (n_14623, out_fifo_read_pointer[0], wc1056);
  not gc1056 (wc1056, out_fifo_write_pointer[0]);
  or g41606 (n_14624, wc1057, out_fifo_write_pointer[0]);
  not gc1057 (wc1057, out_fifo_read_pointer[0]);
  or g41607 (n_14625, out_fifo_read_pointer[2], wc1058);
  not gc1058 (wc1058, out_fifo_write_pointer[2]);
  or g41608 (n_14626, wc1059, out_fifo_write_pointer[2]);
  not gc1059 (wc1059, out_fifo_read_pointer[2]);
  or g41609 (n_20909, wc1060, out_fifo_write_pointer[1]);
  not gc1060 (wc1060, out_fifo_read_pointer[1]);
  or g41610 (n_20910, out_fifo_read_pointer[1], wc1061);
  not gc1061 (wc1061, out_fifo_write_pointer[1]);
  nand g41611 (n_14622, n_20909, n_20910);
  or g41612 (n_12733, wc1062, out_fifo_read_pointer[1]);
  not gc1062 (wc1062, out_fifo_read_pointer[0]);
  or g41613 (n_12734, out_fifo_read_pointer[0], wc1063);
  not gc1063 (wc1063, out_fifo_read_pointer[1]);
  nand g41614 (n_13808, data_stack_pointer[2], rst_n);
  or g41615 (n_13816, data_stack_pointer[0], wc1064);
  not gc1064 (wc1064, rst_n);
  or g41616 (n_14635, sh_reg_out_bit_counter[1],
       sh_reg_out_bit_counter[2]);
  nand g41617 (n_14658, sh_reg_out_bit_counter[0],
       sh_reg_out_bit_counter[1]);
  nand g41618 (n_14648, sh_bit_cnt[0], enable_n);
  or g41619 (n_15633, data_stack_pointer[3], wc1065);
  not gc1065 (wc1065, rst_n);
  or g41620 (n_37, data_stack_pointer[2], data_stack_pointer[3]);
  and g41621 (n_20868, n_14583, wc1066);
  not gc1066 (wc1066, n_11);
  and g41622 (n_20877, wc1067, sh_reg_out[24]);
  not gc1067 (wc1067, n_11);
  and g41623 (n_20878, wc1068, sh_reg_out[23]);
  not gc1068 (wc1068, n_11);
  and g41624 (n_20879, wc1069, sh_reg_out[22]);
  not gc1069 (wc1069, n_11);
  and g41625 (n_20880, wc1070, sh_reg_out[21]);
  not gc1070 (wc1070, n_11);
  and g41626 (n_20881, wc1071, sh_reg_out[8]);
  not gc1071 (wc1071, n_11);
  and g41627 (n_20884, wc1072, sh_reg_out[18]);
  not gc1072 (wc1072, n_11);
  and g41628 (n_20885, wc1073, sh_reg_out[25]);
  not gc1073 (wc1073, n_11);
  and g41629 (n_20886, wc1074, sh_reg_out[26]);
  not gc1074 (wc1074, n_11);
  or g41633 (n_4207, wc1075, n_4175);
  not gc1075 (wc1075, n_14301);
  or g41634 (n_4239, wc1076, n_4207);
  not gc1076 (wc1076, n_14267);
  or g41635 (n_4646, wc1077, n_14480);
  not gc1077 (wc1077, n_3649);
  CDN_flop \out_fifo_read_pointer_reg[0] (.clk (clk), .d (n_5023),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[0]));
  CDN_flop \out_fifo_read_pointer_reg[1] (.clk (clk), .d (n_5027),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[1]));
  CDN_flop \out_fifo_read_pointer_reg[2] (.clk (clk), .d (n_5031),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[2]));
  CDN_flop \out_fifo_reg[0][0][0] (.clk (clk), .d (n_5715), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [0]));
  CDN_flop \out_fifo_reg[0][0][1] (.clk (clk), .d (n_5035), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [1]));
  CDN_flop \out_fifo_reg[0][0][2] (.clk (clk), .d (n_5039), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [2]));
  CDN_flop \out_fifo_reg[0][0][3] (.clk (clk), .d (n_5043), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [3]));
  CDN_flop \out_fifo_reg[0][0][4] (.clk (clk), .d (n_5047), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [4]));
  CDN_flop \out_fifo_reg[0][0][5] (.clk (clk), .d (n_5051), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [5]));
  CDN_flop \out_fifo_reg[0][0][6] (.clk (clk), .d (n_5055), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [6]));
  CDN_flop \out_fifo_reg[0][0][7] (.clk (clk), .d (n_5059), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [7]));
  CDN_flop \out_fifo_reg[0][0][8] (.clk (clk), .d (n_5063), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [8]));
  CDN_flop \out_fifo_reg[0][1][0] (.clk (clk), .d (n_5747), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [0]));
  CDN_flop \out_fifo_reg[0][1][1] (.clk (clk), .d (n_5067), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [1]));
  CDN_flop \out_fifo_reg[0][1][2] (.clk (clk), .d (n_5071), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [2]));
  CDN_flop \out_fifo_reg[0][1][3] (.clk (clk), .d (n_5075), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [3]));
  CDN_flop \out_fifo_reg[0][1][4] (.clk (clk), .d (n_5079), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [4]));
  CDN_flop \out_fifo_reg[0][1][5] (.clk (clk), .d (n_5083), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [5]));
  CDN_flop \out_fifo_reg[0][1][6] (.clk (clk), .d (n_5087), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [6]));
  CDN_flop \out_fifo_reg[0][1][7] (.clk (clk), .d (n_5091), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [7]));
  CDN_flop \out_fifo_reg[0][1][8] (.clk (clk), .d (n_5095), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [8]));
  CDN_flop \out_fifo_reg[0][2][0] (.clk (clk), .d (n_5779), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [0]));
  CDN_flop \out_fifo_reg[0][2][1] (.clk (clk), .d (n_5099), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [1]));
  CDN_flop \out_fifo_reg[0][2][8] (.clk (clk), .d (n_5103), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [8]));
  CDN_flop \out_fifo_reg[0][2][9] (.clk (clk), .d (1'b1), .sena
       (n_887), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (\out_fifo[0][2] [9]));
  CDN_flop \out_fifo_reg[1][0][0] (.clk (clk), .d (n_5719), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [0]));
  CDN_flop \out_fifo_reg[1][0][1] (.clk (clk), .d (n_5107), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [1]));
  CDN_flop \out_fifo_reg[1][0][2] (.clk (clk), .d (n_5111), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [2]));
  CDN_flop \out_fifo_reg[1][0][3] (.clk (clk), .d (n_5115), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [3]));
  CDN_flop \out_fifo_reg[1][0][4] (.clk (clk), .d (n_5119), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [4]));
  CDN_flop \out_fifo_reg[1][0][5] (.clk (clk), .d (n_5123), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [5]));
  CDN_flop \out_fifo_reg[1][0][6] (.clk (clk), .d (n_5127), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [6]));
  CDN_flop \out_fifo_reg[1][0][7] (.clk (clk), .d (n_5131), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [7]));
  CDN_flop \out_fifo_reg[1][0][8] (.clk (clk), .d (n_5135), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [8]));
  CDN_flop \out_fifo_reg[1][1][0] (.clk (clk), .d (n_5751), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [0]));
  CDN_flop \out_fifo_reg[1][1][1] (.clk (clk), .d (n_5139), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [1]));
  CDN_flop \out_fifo_reg[1][1][2] (.clk (clk), .d (n_5143), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [2]));
  CDN_flop \out_fifo_reg[1][1][3] (.clk (clk), .d (n_5147), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [3]));
  CDN_flop \out_fifo_reg[1][1][4] (.clk (clk), .d (n_5151), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [4]));
  CDN_flop \out_fifo_reg[1][1][5] (.clk (clk), .d (n_5155), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [5]));
  CDN_flop \out_fifo_reg[1][1][6] (.clk (clk), .d (n_5159), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [6]));
  CDN_flop \out_fifo_reg[1][1][7] (.clk (clk), .d (n_5163), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [7]));
  CDN_flop \out_fifo_reg[1][1][8] (.clk (clk), .d (n_5167), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [8]));
  CDN_flop \out_fifo_reg[1][2][0] (.clk (clk), .d (n_5783), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [0]));
  CDN_flop \out_fifo_reg[1][2][1] (.clk (clk), .d (n_5171), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [1]));
  CDN_flop \out_fifo_reg[1][2][8] (.clk (clk), .d (n_5175), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [8]));
  CDN_flop \out_fifo_reg[1][2][9] (.clk (clk), .d (1'b1), .sena
       (n_877), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (\out_fifo[1][2] [9]));
  CDN_flop \out_fifo_reg[2][0][0] (.clk (clk), .d (n_5723), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [0]));
  CDN_flop \out_fifo_reg[2][0][1] (.clk (clk), .d (n_5179), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [1]));
  CDN_flop \out_fifo_reg[2][0][2] (.clk (clk), .d (n_5183), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [2]));
  CDN_flop \out_fifo_reg[2][0][3] (.clk (clk), .d (n_5187), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [3]));
  CDN_flop \out_fifo_reg[2][0][4] (.clk (clk), .d (n_5191), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [4]));
  CDN_flop \out_fifo_reg[2][0][5] (.clk (clk), .d (n_5195), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [5]));
  CDN_flop \out_fifo_reg[2][0][6] (.clk (clk), .d (n_5199), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [6]));
  CDN_flop \out_fifo_reg[2][0][7] (.clk (clk), .d (n_5203), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [7]));
  CDN_flop \out_fifo_reg[2][0][8] (.clk (clk), .d (n_5207), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [8]));
  CDN_flop \out_fifo_reg[2][1][0] (.clk (clk), .d (n_5755), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [0]));
  CDN_flop \out_fifo_reg[2][1][1] (.clk (clk), .d (n_5211), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [1]));
  CDN_flop \out_fifo_reg[2][1][2] (.clk (clk), .d (n_5215), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [2]));
  CDN_flop \out_fifo_reg[2][1][3] (.clk (clk), .d (n_5219), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [3]));
  CDN_flop \out_fifo_reg[2][1][4] (.clk (clk), .d (n_5223), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [4]));
  CDN_flop \out_fifo_reg[2][1][5] (.clk (clk), .d (n_5227), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [5]));
  CDN_flop \out_fifo_reg[2][1][6] (.clk (clk), .d (n_5231), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [6]));
  CDN_flop \out_fifo_reg[2][1][7] (.clk (clk), .d (n_5235), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [7]));
  CDN_flop \out_fifo_reg[2][1][8] (.clk (clk), .d (n_5239), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [8]));
  CDN_flop \out_fifo_reg[2][2][0] (.clk (clk), .d (n_5787), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [0]));
  CDN_flop \out_fifo_reg[2][2][1] (.clk (clk), .d (n_5243), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [1]));
  CDN_flop \out_fifo_reg[2][2][8] (.clk (clk), .d (n_5247), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [8]));
  CDN_flop \out_fifo_reg[2][2][9] (.clk (clk), .d (1'b1), .sena
       (n_867), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (\out_fifo[2][2] [9]));
  CDN_flop \out_fifo_reg[3][0][0] (.clk (clk), .d (n_5727), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [0]));
  CDN_flop \out_fifo_reg[3][0][1] (.clk (clk), .d (n_5251), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [1]));
  CDN_flop \out_fifo_reg[3][0][2] (.clk (clk), .d (n_5255), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [2]));
  CDN_flop \out_fifo_reg[3][0][3] (.clk (clk), .d (n_5259), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [3]));
  CDN_flop \out_fifo_reg[3][0][4] (.clk (clk), .d (n_5263), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [4]));
  CDN_flop \out_fifo_reg[3][0][5] (.clk (clk), .d (n_5267), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [5]));
  CDN_flop \out_fifo_reg[3][0][6] (.clk (clk), .d (n_5271), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [6]));
  CDN_flop \out_fifo_reg[3][0][7] (.clk (clk), .d (n_5275), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [7]));
  CDN_flop \out_fifo_reg[3][0][8] (.clk (clk), .d (n_5279), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [8]));
  CDN_flop \out_fifo_reg[3][1][0] (.clk (clk), .d (n_5759), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [0]));
  CDN_flop \out_fifo_reg[3][1][1] (.clk (clk), .d (n_5283), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [1]));
  CDN_flop \out_fifo_reg[3][1][2] (.clk (clk), .d (n_5287), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [2]));
  CDN_flop \out_fifo_reg[3][1][3] (.clk (clk), .d (n_5291), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [3]));
  CDN_flop \out_fifo_reg[3][1][4] (.clk (clk), .d (n_5295), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [4]));
  CDN_flop \out_fifo_reg[3][1][5] (.clk (clk), .d (n_5299), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [5]));
  CDN_flop \out_fifo_reg[3][1][6] (.clk (clk), .d (n_5303), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [6]));
  CDN_flop \out_fifo_reg[3][1][7] (.clk (clk), .d (n_5307), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [7]));
  CDN_flop \out_fifo_reg[3][1][8] (.clk (clk), .d (n_5311), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [8]));
  CDN_flop \out_fifo_reg[3][2][0] (.clk (clk), .d (n_5791), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [0]));
  CDN_flop \out_fifo_reg[3][2][1] (.clk (clk), .d (n_5315), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [1]));
  CDN_flop \out_fifo_reg[3][2][8] (.clk (clk), .d (n_5319), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [8]));
  CDN_flop \out_fifo_reg[3][2][9] (.clk (clk), .d (1'b1), .sena
       (n_20862), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd
       (1'b0), .q (\out_fifo[3][2] [9]));
  CDN_flop \out_fifo_reg[4][0][0] (.clk (clk), .d (n_5731), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [0]));
  CDN_flop \out_fifo_reg[4][0][1] (.clk (clk), .d (n_5323), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [1]));
  CDN_flop \out_fifo_reg[4][0][2] (.clk (clk), .d (n_5327), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [2]));
  CDN_flop \out_fifo_reg[4][0][3] (.clk (clk), .d (n_5331), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [3]));
  CDN_flop \out_fifo_reg[4][0][4] (.clk (clk), .d (n_5335), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [4]));
  CDN_flop \out_fifo_reg[4][0][5] (.clk (clk), .d (n_5339), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [5]));
  CDN_flop \out_fifo_reg[4][0][6] (.clk (clk), .d (n_5343), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [6]));
  CDN_flop \out_fifo_reg[4][0][7] (.clk (clk), .d (n_5347), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [7]));
  CDN_flop \out_fifo_reg[4][0][8] (.clk (clk), .d (n_5351), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [8]));
  CDN_flop \out_fifo_reg[4][1][0] (.clk (clk), .d (n_5763), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [0]));
  CDN_flop \out_fifo_reg[4][1][1] (.clk (clk), .d (n_5355), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [1]));
  CDN_flop \out_fifo_reg[4][1][2] (.clk (clk), .d (n_5359), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [2]));
  CDN_flop \out_fifo_reg[4][1][3] (.clk (clk), .d (n_5363), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [3]));
  CDN_flop \out_fifo_reg[4][1][4] (.clk (clk), .d (n_5367), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [4]));
  CDN_flop \out_fifo_reg[4][1][5] (.clk (clk), .d (n_5371), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [5]));
  CDN_flop \out_fifo_reg[4][1][6] (.clk (clk), .d (n_5375), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [6]));
  CDN_flop \out_fifo_reg[4][1][7] (.clk (clk), .d (n_5379), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [7]));
  CDN_flop \out_fifo_reg[4][1][8] (.clk (clk), .d (n_5383), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [8]));
  CDN_flop \out_fifo_reg[4][2][0] (.clk (clk), .d (n_5795), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [0]));
  CDN_flop \out_fifo_reg[4][2][1] (.clk (clk), .d (n_5387), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [1]));
  CDN_flop \out_fifo_reg[4][2][8] (.clk (clk), .d (n_5391), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [8]));
  CDN_flop \out_fifo_reg[4][2][9] (.clk (clk), .d (1'b1), .sena
       (n_847), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (\out_fifo[4][2] [9]));
  CDN_flop \out_fifo_reg[5][0][0] (.clk (clk), .d (n_5735), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [0]));
  CDN_flop \out_fifo_reg[5][0][1] (.clk (clk), .d (n_5395), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [1]));
  CDN_flop \out_fifo_reg[5][0][2] (.clk (clk), .d (n_5399), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [2]));
  CDN_flop \out_fifo_reg[5][0][3] (.clk (clk), .d (n_5403), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [3]));
  CDN_flop \out_fifo_reg[5][0][4] (.clk (clk), .d (n_5407), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [4]));
  CDN_flop \out_fifo_reg[5][0][5] (.clk (clk), .d (n_5411), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [5]));
  CDN_flop \out_fifo_reg[5][0][6] (.clk (clk), .d (n_5415), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [6]));
  CDN_flop \out_fifo_reg[5][0][7] (.clk (clk), .d (n_5419), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [7]));
  CDN_flop \out_fifo_reg[5][0][8] (.clk (clk), .d (n_5423), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [8]));
  CDN_flop \out_fifo_reg[5][1][0] (.clk (clk), .d (n_5767), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [0]));
  CDN_flop \out_fifo_reg[5][1][1] (.clk (clk), .d (n_5427), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [1]));
  CDN_flop \out_fifo_reg[5][1][2] (.clk (clk), .d (n_5431), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [2]));
  CDN_flop \out_fifo_reg[5][1][3] (.clk (clk), .d (n_5435), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [3]));
  CDN_flop \out_fifo_reg[5][1][4] (.clk (clk), .d (n_5439), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [4]));
  CDN_flop \out_fifo_reg[5][1][5] (.clk (clk), .d (n_5443), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [5]));
  CDN_flop \out_fifo_reg[5][1][6] (.clk (clk), .d (n_5447), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [6]));
  CDN_flop \out_fifo_reg[5][1][7] (.clk (clk), .d (n_5451), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [7]));
  CDN_flop \out_fifo_reg[5][1][8] (.clk (clk), .d (n_5455), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [8]));
  CDN_flop \out_fifo_reg[5][2][0] (.clk (clk), .d (n_5799), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [0]));
  CDN_flop \out_fifo_reg[5][2][1] (.clk (clk), .d (n_5459), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [1]));
  CDN_flop \out_fifo_reg[5][2][8] (.clk (clk), .d (n_5463), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [8]));
  CDN_flop \out_fifo_reg[5][2][9] (.clk (clk), .d (1'b1), .sena
       (n_837), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (\out_fifo[5][2] [9]));
  CDN_flop \out_fifo_reg[6][0][0] (.clk (clk), .d (n_5739), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [0]));
  CDN_flop \out_fifo_reg[6][0][1] (.clk (clk), .d (n_5467), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [1]));
  CDN_flop \out_fifo_reg[6][0][2] (.clk (clk), .d (n_5471), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [2]));
  CDN_flop \out_fifo_reg[6][0][3] (.clk (clk), .d (n_5475), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [3]));
  CDN_flop \out_fifo_reg[6][0][4] (.clk (clk), .d (n_5479), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [4]));
  CDN_flop \out_fifo_reg[6][0][5] (.clk (clk), .d (n_5483), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [5]));
  CDN_flop \out_fifo_reg[6][0][6] (.clk (clk), .d (n_5487), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [6]));
  CDN_flop \out_fifo_reg[6][0][7] (.clk (clk), .d (n_5491), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [7]));
  CDN_flop \out_fifo_reg[6][0][8] (.clk (clk), .d (n_5495), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [8]));
  CDN_flop \out_fifo_reg[6][1][0] (.clk (clk), .d (n_5771), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [0]));
  CDN_flop \out_fifo_reg[6][1][1] (.clk (clk), .d (n_5499), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [1]));
  CDN_flop \out_fifo_reg[6][1][2] (.clk (clk), .d (n_5503), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [2]));
  CDN_flop \out_fifo_reg[6][1][3] (.clk (clk), .d (n_5507), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [3]));
  CDN_flop \out_fifo_reg[6][1][4] (.clk (clk), .d (n_5511), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [4]));
  CDN_flop \out_fifo_reg[6][1][5] (.clk (clk), .d (n_5515), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [5]));
  CDN_flop \out_fifo_reg[6][1][6] (.clk (clk), .d (n_5519), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [6]));
  CDN_flop \out_fifo_reg[6][1][7] (.clk (clk), .d (n_5523), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [7]));
  CDN_flop \out_fifo_reg[6][1][8] (.clk (clk), .d (n_5527), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [8]));
  CDN_flop \out_fifo_reg[6][2][0] (.clk (clk), .d (n_5803), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [0]));
  CDN_flop \out_fifo_reg[6][2][1] (.clk (clk), .d (n_5531), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [1]));
  CDN_flop \out_fifo_reg[6][2][8] (.clk (clk), .d (n_5535), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [8]));
  CDN_flop \out_fifo_reg[6][2][9] (.clk (clk), .d (1'b1), .sena
       (n_827), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (\out_fifo[6][2] [9]));
  CDN_flop \out_fifo_reg[7][0][0] (.clk (clk), .d (n_5743), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [0]));
  CDN_flop \out_fifo_reg[7][0][1] (.clk (clk), .d (n_5539), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [1]));
  CDN_flop \out_fifo_reg[7][0][2] (.clk (clk), .d (n_5543), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [2]));
  CDN_flop \out_fifo_reg[7][0][3] (.clk (clk), .d (n_5547), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [3]));
  CDN_flop \out_fifo_reg[7][0][4] (.clk (clk), .d (n_5551), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [4]));
  CDN_flop \out_fifo_reg[7][0][5] (.clk (clk), .d (n_5555), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [5]));
  CDN_flop \out_fifo_reg[7][0][6] (.clk (clk), .d (n_5559), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [6]));
  CDN_flop \out_fifo_reg[7][0][7] (.clk (clk), .d (n_5563), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [7]));
  CDN_flop \out_fifo_reg[7][0][8] (.clk (clk), .d (n_5567), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [8]));
  CDN_flop \out_fifo_reg[7][1][0] (.clk (clk), .d (n_5775), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [0]));
  CDN_flop \out_fifo_reg[7][1][1] (.clk (clk), .d (n_5571), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [1]));
  CDN_flop \out_fifo_reg[7][1][2] (.clk (clk), .d (n_5575), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [2]));
  CDN_flop \out_fifo_reg[7][1][3] (.clk (clk), .d (n_5579), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [3]));
  CDN_flop \out_fifo_reg[7][1][4] (.clk (clk), .d (n_5583), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [4]));
  CDN_flop \out_fifo_reg[7][1][5] (.clk (clk), .d (n_5587), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [5]));
  CDN_flop \out_fifo_reg[7][1][6] (.clk (clk), .d (n_5591), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [6]));
  CDN_flop \out_fifo_reg[7][1][7] (.clk (clk), .d (n_5595), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [7]));
  CDN_flop \out_fifo_reg[7][1][8] (.clk (clk), .d (n_5599), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [8]));
  CDN_flop \out_fifo_reg[7][2][0] (.clk (clk), .d (n_5807), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [0]));
  CDN_flop \out_fifo_reg[7][2][1] (.clk (clk), .d (n_5603), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [1]));
  CDN_flop \out_fifo_reg[7][2][8] (.clk (clk), .d (n_5607), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [8]));
  CDN_flop \out_fifo_reg[7][2][9] (.clk (clk), .d (1'b1), .sena
       (n_20863), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd
       (1'b0), .q (\out_fifo[7][2] [9]));
  CDN_flop \out_fifo_write_pointer_reg[0] (.clk (clk), .d (n_5611),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[0]));
  CDN_flop \out_fifo_write_pointer_reg[1] (.clk (clk), .d (n_5615),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[1]));
  CDN_flop \out_fifo_write_pointer_reg[2] (.clk (clk), .d (n_5619),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[2]));
  CDN_flop \sh_bit_cnt_reg[0] (.clk (clk), .d (n_5622), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[0]));
  CDN_flop \sh_bit_cnt_reg[1] (.clk (clk), .d (n_5625), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[1]));
  CDN_flop \sh_bit_cnt_reg[2] (.clk (clk), .d (n_5628), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[2]));
  CDN_flop \sh_bit_cnt_reg[3] (.clk (clk), .d (n_5631), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[3]));
  CDN_flop \sh_reg_in_reg[0] (.clk (clk), .d (din), .sena (n_523),
       .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0), .q
       (sh_reg_in[0]));
  CDN_flop \sh_reg_in_reg[1] (.clk (clk), .d (sh_reg_in[0]), .sena
       (n_523), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (sh_reg_in[1]));
  CDN_flop \sh_reg_in_reg[2] (.clk (clk), .d (sh_reg_in[1]), .sena
       (n_523), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (sh_reg_in[2]));
  CDN_flop \sh_reg_in_reg[3] (.clk (clk), .d (sh_reg_in[2]), .sena
       (n_523), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (sh_reg_in[3]));
  CDN_flop \sh_reg_in_reg[4] (.clk (clk), .d (sh_reg_in[3]), .sena
       (n_523), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (sh_reg_in[4]));
  CDN_flop \sh_reg_in_reg[5] (.clk (clk), .d (sh_reg_in[4]), .sena
       (n_523), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (sh_reg_in[5]));
  CDN_flop \sh_reg_in_reg[6] (.clk (clk), .d (sh_reg_in[5]), .sena
       (n_523), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (sh_reg_in[6]));
  CDN_flop \sh_reg_in_reg[7] (.clk (clk), .d (sh_reg_in[6]), .sena
       (n_523), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (sh_reg_in[7]));
  CDN_flop \sh_reg_in_reg[8] (.clk (clk), .d (sh_reg_in[7]), .sena
       (n_523), .aclr (1'b0), .apre (1'b0), .srl (n_521), .srd (1'b0),
       .q (sh_reg_in[8]));
  CDN_flop \sh_reg_out_bit_counter_reg[0] (.clk (clk), .d (n_5635),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[0]));
  CDN_flop \sh_reg_out_bit_counter_reg[1] (.clk (clk), .d (n_20868),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[1]));
  CDN_flop \sh_reg_out_bit_counter_reg[2] (.clk (clk), .d (n_5643),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[2]));
  CDN_flop \sh_reg_out_bit_counter_reg[3] (.clk (clk), .d (n_5647),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[3]));
  CDN_flop \sh_reg_out_bit_counter_reg[4] (.clk (clk), .d (n_5651),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[4]));
  CDN_flop \sh_reg_out_reg[0] (.clk (clk), .d (n_5653), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[0]));
  CDN_flop \sh_reg_out_reg[1] (.clk (clk), .d (n_5655), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[1]));
  CDN_flop \sh_reg_out_reg[2] (.clk (clk), .d (n_5657), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[2]));
  CDN_flop \sh_reg_out_reg[3] (.clk (clk), .d (n_5659), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[3]));
  CDN_flop \sh_reg_out_reg[4] (.clk (clk), .d (n_5661), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[4]));
  CDN_flop \sh_reg_out_reg[5] (.clk (clk), .d (n_5663), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[5]));
  CDN_flop \sh_reg_out_reg[6] (.clk (clk), .d (n_5665), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[6]));
  CDN_flop \sh_reg_out_reg[7] (.clk (clk), .d (n_5667), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[7]));
  CDN_flop \sh_reg_out_reg[8] (.clk (clk), .d (n_5669), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[8]));
  CDN_flop \sh_reg_out_reg[9] (.clk (clk), .d (n_20881), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[9]));
  CDN_flop \sh_reg_out_reg[10] (.clk (clk), .d (n_5673), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[10]));
  CDN_flop \sh_reg_out_reg[11] (.clk (clk), .d (n_5675), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[11]));
  CDN_flop \sh_reg_out_reg[12] (.clk (clk), .d (n_5677), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[12]));
  CDN_flop \sh_reg_out_reg[13] (.clk (clk), .d (n_5679), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[13]));
  CDN_flop \sh_reg_out_reg[14] (.clk (clk), .d (n_5681), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[14]));
  CDN_flop \sh_reg_out_reg[15] (.clk (clk), .d (n_5683), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[15]));
  CDN_flop \sh_reg_out_reg[16] (.clk (clk), .d (n_5685), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[16]));
  CDN_flop \sh_reg_out_reg[17] (.clk (clk), .d (n_5687), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[17]));
  CDN_flop \sh_reg_out_reg[18] (.clk (clk), .d (n_5689), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[18]));
  CDN_flop \sh_reg_out_reg[19] (.clk (clk), .d (n_20884), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[19]));
  CDN_flop \sh_reg_out_reg[20] (.clk (clk), .d (n_5693), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[20]));
  CDN_flop \sh_reg_out_reg[21] (.clk (clk), .d (n_5695), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[21]));
  CDN_flop \sh_reg_out_reg[22] (.clk (clk), .d (n_20880), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[22]));
  CDN_flop \sh_reg_out_reg[23] (.clk (clk), .d (n_20879), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[23]));
  CDN_flop \sh_reg_out_reg[24] (.clk (clk), .d (n_20878), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[24]));
  CDN_flop \sh_reg_out_reg[25] (.clk (clk), .d (n_20877), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[25]));
  CDN_flop \sh_reg_out_reg[26] (.clk (clk), .d (n_20885), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[26]));
  CDN_flop \sh_reg_out_reg[27] (.clk (clk), .d (n_20886), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[27]));
  CDN_flop \sh_reg_out_reg[28] (.clk (clk), .d (n_5709), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[28]));
  CDN_flop \sh_reg_out_reg[29] (.clk (clk), .d (n_5711), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (dout));
endmodule

`ifdef RC_CDN_GENERIC_GATE
`else
module CDN_flop(clk, d, sena, aclr, apre, srl, srd, q);
  input clk, d, sena, aclr, apre, srl, srd;
  output q;
  wire clk, d, sena, aclr, apre, srl, srd;
  wire q;
  reg  qi;
  assign #1 q = qi;
  always 
    @(posedge clk or posedge apre or posedge aclr) 
      if (aclr) 
        qi <= 0;
      else if (apre) 
          qi <= 1;
        else if (srl) 
            qi <= srd;
          else begin
            if (sena) 
              qi <= d;
          end
  initial 
    qi <= 1'b0;
endmodule
`endif
