/*
 Copyright 2013 Ray Salemi

 Licensed under the Apache License, Version 2.0 (the "License");
 you may not use this file except in compliance with the License.
 You may obtain a copy of the License at

 http://www.apache.org/licenses/LICENSE-2.0

 Unless required by applicable law or agreed to in writing, software
 distributed under the License is distributed on an "AS IS" BASIS,
 WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 See the License for the specific language governing permissions and
 limitations under the License.
 */
class vdic_dut_reset_sequence extends uvm_sequence #(vdic_dut_sequence_item);
    `uvm_object_utils(vdic_dut_reset_sequence)

//------------------------------------------------------------------------------
// local variables
//------------------------------------------------------------------------------

// Not necessary: req is inherited
//    sequence_item req;

//------------------------------------------------------------------------------
// constructor
//------------------------------------------------------------------------------

    function new(string name = "reset");
        super.new(name);
    endfunction : new
    
//------------------------------------------------------------------------------
// the sequence body
//------------------------------------------------------------------------------

    task body();
        `uvm_info("SEQ_RESET", "", UVM_MEDIUM)
        `uvm_do_with(req, {state == RESET;} )
    endtask : body
    
    
endclass : vdic_dut_reset_sequence












