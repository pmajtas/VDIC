/******************************************************************************
 * (C) Copyright 2022 AGH UST All Rights Reserved
 ******************************************************************************
 * MODULE NAME: vdic_dut_2022
 * VERSION:     1.0
 * DATE:        21-10-2022
 *
 * ABSTRACT:   DUT module for VDIC 2022 labs.
 *              The DUT is RPN calculator type. The arguments are sent first,
 *              than the operator/command.
 *******************************************************************************
 * INPUTS
 *    clk      - posedge active clock, always running
 *    rst_n    - synchronous reset active low
 *    din      - serial data input
 *    enable_n - chip enable, active low;

 * OUTPUTS
 *    dout       - serial data output
 *    dout_valid - valid flag for serial data output, active high
 *
 *******************************************************************************

 The clock is always active.
 The DUT operates on the posedge of the clock.
 The DUT receives the data when enable_n is active.

 --------------------------------------------------------------------------------
 --- Input data
 --------------------------------------------------------------------------------

 The input data is send serially in WORDs.

 The WORD is always 10 bit long. MSB is sent first.
 The WORD sent to the DUT is either DATA type or CONTROL type.

 DATA = 0bbbbbbbbp
 where:
 - b = 0 or 1, PAYLOAD bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 CONTROL = 1bbbbbbbbp
 where:
 - b = 0 or 1, COMMAND bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 The COMMAND can be:
 00000000 - CMD_NOP, do nothing, remove the data (reset data stack)
 00000001 - CMD_AND, logic AND of the last two arguments
 00000010 - CMD_OR, logic OR of the arguments
 00000011 - CMD_XOR, logic XOR of the arguments
 00010000 - CMD_ADD, add the arguments
 00100000 - CMD_SUB, subtract other arguments from the first one

 --------------------------------------------------------------------------------
 --- Output data
 --------------------------------------------------------------------------------

 The DUT responds to each CONTROL word, sending 3 WORDS:
 STATUS, DATA, DATA

 STATUS = 1bbbbbbbbp
 where bbbbbbbb is one of:

 00000000 - S_NO_ERROR - data correctly processed
 00000001 - S_MISSING_DATA - missing input data
 00000010 - S_DATA_STACK_OVERFLOW - maximum number of arguments exceeded
 00000100 - S_OUTPUT_FIFO_OVERFLOW - result dropped not possible to process
 00100000 - S_DATA_PARITY_ERROR - input data or command parity error
 01000000 - S_COMMAND_PARITY_ERROR - input data or command parity error
 10000000 - S_INVALID_COMMAND - unknown command detected

 DATA is defined as in the input.
 PAYLOAD of the DATA is 00000000 if the data was NOT processed correctly.

 *******************************************************************************
 * IMPLEMENTATION STATUS
 *******************************************************************************
 *  <Feature>                        <Is implemented>
 *    command CMD_NOP                    NO
 *    command CMD_AND                   YES
 *    command CMD_OR                     NO
 *    command CMD_XOR                    NO
 *    command CMD_ADD                   YES
 *    command CMD_SUB                    NO
 *    status S_NO_ERROR                 YES
 *    status S_MISSING_DATA              NO
 *    status S_DATA_STACK_OVERFLOW       NO
 *    status S_OUTPUT_FIFO_OVERFLOW      NO
 *    status S_DATA_PARITY_ERROR         NO
 *    status S_COMMAND_PARITY_ERROR      NO
 *    status S_INVALID_COMMAND          YES
 *******************************************************************************
 */

// Generated by Cadence Genus(TM) Synthesis Solution 19.15-s090_1
// Generated on: Oct 20 2022 12:35:05 CEST (Oct 20 2022 10:35:05 UTC)

// Verification Directory ./LEC 

module vdic_dut_2022(clk, rst_n, enable_n, din, dout, dout_valid);
  input clk, rst_n, enable_n, din;
  output dout, dout_valid;
  wire clk, rst_n, enable_n, din;
  wire dout, dout_valid;
  wire [7:0] \data_stack_mem[0] ;
  wire [7:0] \data_stack_mem[1] ;
  wire [7:0] \data_stack_mem[2] ;
  wire [7:0] \data_stack_mem[3] ;
  wire [7:0] \data_stack_mem[4] ;
  wire [7:0] \data_stack_mem[5] ;
  wire [7:0] \data_stack_mem[6] ;
  wire [7:0] \data_stack_mem[7] ;
  wire [7:0] \data_stack_mem[8] ;
  wire [3:0] data_stack_pointer;
  wire [2:0] out_fifo_write_pointer;
  wire [3:0] sh_bit_cnt;
  wire [4:0] sh_reg_out_bit_counter;
  wire [2:0] out_fifo_read_pointer;
  wire [9:0] sh_reg_in;
  wire [9:0] \out_fifo[0][1] ;
  wire [9:0] \out_fifo[4][0] ;
  wire [9:0] \out_fifo[0][0] ;
  wire [9:0] \out_fifo[4][1] ;
  wire [9:0] \out_fifo[0][2] ;
  wire [9:0] \out_fifo[4][2] ;
  wire [9:0] \out_fifo[2][0] ;
  wire [9:0] \out_fifo[1][0] ;
  wire [9:0] \out_fifo[3][0] ;
  wire [9:0] \out_fifo[5][0] ;
  wire [9:0] \out_fifo[6][0] ;
  wire [9:0] \out_fifo[7][0] ;
  wire [9:0] \out_fifo[2][2] ;
  wire [9:0] \out_fifo[1][2] ;
  wire [9:0] \out_fifo[3][2] ;
  wire [9:0] \out_fifo[5][2] ;
  wire [9:0] \out_fifo[6][2] ;
  wire [9:0] \out_fifo[7][2] ;
  wire [9:0] \out_fifo[2][1] ;
  wire [9:0] \out_fifo[1][1] ;
  wire [9:0] \out_fifo[3][1] ;
  wire [9:0] \out_fifo[5][1] ;
  wire [9:0] \out_fifo[6][1] ;
  wire [9:0] \out_fifo[7][1] ;
  wire [29:0] sh_reg_out;
  wire n_11453, n_11454, n_11455, n_11456, n_11457, n_11462, n_11463,
       n_11468;
  wire n_11469, n_11470, n_11475, n_11476, n_11477, n_11478, n_11479,
       n_11480;
  wire n_11481, n_11482, n_11483, n_11484, n_11485, n_11486, n_11487,
       n_11488;
  wire n_11489, n_11490, n_11491, n_11492, n_11493, n_11494, n_11495,
       n_11496;
  wire n_11497, n_11498, n_11500, n_11501, n_11502, n_11503, n_11504,
       n_11505;
  wire n_11506, n_11507, n_11508, n_11509, n_11510, n_11511, n_11512,
       n_11513;
  wire n_11514, n_11515, n_11516, n_11517, n_11518, n_11519, n_11520,
       n_11521;
  wire n_11522, n_11523, n_11524, n_11525, n_11526, n_11527, n_11528,
       n_11529;
  wire n_11530, n_11531, n_11532, n_11533, n_11534, n_11535, n_11536,
       n_11537;
  wire n_11538, n_11539, n_11540, n_11541, n_11542, n_11543, n_11544,
       n_11545;
  wire n_11546, n_11547, n_11548, n_11549, n_11550, n_11551, n_11552,
       n_11553;
  wire n_11554, n_11555, n_11556, n_11557, n_11558, n_11559, n_11560,
       n_11561;
  wire n_11562, n_11563, n_11564, n_11565, n_11566, n_11567, n_11568,
       n_11569;
  wire n_11570, n_11571, n_11572, n_11573, n_11574, n_11575, n_11576,
       n_11577;
  wire n_11578, n_11579, n_11580, n_11581, n_11582, n_11583, n_11584,
       n_11585;
  wire n_11586, n_11587, n_11588, n_11589, n_11590, n_11591, n_11592,
       n_11593;
  wire n_11594, n_11595, n_11596, n_11597, n_11598, n_11599, n_11600,
       n_11601;
  wire n_11602, n_11603, n_11604, n_11605, n_11606, n_11607, n_11608,
       n_11609;
  wire n_11610, n_11611, n_11612, n_11613, n_11614, n_11615, n_11616,
       n_11617;
  wire n_11618, n_11619, n_11621, n_11622, n_11623, n_11624, n_11625,
       n_11626;
  wire n_11627, n_11628, n_11629, n_11630, n_11631, n_11632, n_11633,
       n_11634;
  wire n_11635, n_11636, n_11637, n_11638, n_11639, n_11640, n_11641,
       n_11642;
  wire n_11643, n_11644, n_11645, n_11646, n_11647, n_11648, n_11649,
       n_11650;
  wire n_11651, n_11652, n_11654, n_11655, n_11656, n_11657, n_11658,
       n_11659;
  wire n_11660, n_11661, n_11662, n_11663, n_11664, n_11665, n_11666,
       n_11667;
  wire n_11668, n_11669, n_11670, n_11671, n_11672, n_11673, n_11674,
       n_11675;
  wire n_11676, n_11677, n_11678, n_11679, n_11680, n_11681, n_11682,
       n_11683;
  wire n_11684, n_11685, n_11686, n_11687, n_11688, n_11689, n_11690,
       n_11691;
  wire n_11692, n_11693, n_11694, n_11695, n_11696, n_11697, n_11698,
       n_11699;
  wire n_11700, n_11701, n_11702, n_11703, n_11704, n_11705, n_11706,
       n_11707;
  wire n_11708, n_11709, n_11710, n_11711, n_11712, n_11713, n_11714,
       n_11715;
  wire n_11716, n_11717, n_11718, n_11719, n_11720, n_11721, n_11722,
       n_11723;
  wire n_11724, n_11725, n_11726, n_11727, n_11728, n_11729, n_11730,
       n_11731;
  wire n_11732, n_11733, n_11734, n_11735, n_11736, n_11737, n_11738,
       n_11739;
  wire n_11740, n_11741, n_11742, n_11743, n_11744, n_11745, n_11746,
       n_11747;
  wire n_11748, n_11749, n_11750, n_11751, n_11752, n_11753, n_11754,
       n_11755;
  wire n_11756, n_11757, n_11758, n_11759, n_11760, n_11761, n_11762,
       n_11763;
  wire n_11764, n_11765, n_11766, n_11767, n_11768, n_11769, n_11770,
       n_11771;
  wire n_11772, n_11773, n_11774, n_11775, n_11776, n_11777, n_11778,
       n_11779;
  wire n_11780, n_11781, n_11782, n_11783, n_11784, n_11785, n_11786,
       n_11787;
  wire n_11788, n_11789, n_11790, n_11791, n_11792, n_11793, n_11794,
       n_11795;
  wire n_11796, n_11797, n_11798, n_11799, n_11800, n_11801, n_11802,
       n_11803;
  wire n_11804, n_11805, n_11806, n_11807, n_11808, n_11809, n_11810,
       n_11811;
  wire n_11812, n_11813, n_11815, n_11816, n_11817, n_11818, n_11819,
       n_11820;
  wire n_11821, n_11822, n_11823, n_11824, n_11825, n_11826, n_11827,
       n_11828;
  wire n_11829, n_11830, n_11831, n_11832, n_11833, n_11834, n_11835,
       n_11836;
  wire n_11837, n_11838, n_11839, n_11840, n_11841, n_11842, n_11843,
       n_11844;
  wire n_11845, n_11846, n_11847, n_11848, n_11849, n_11850, n_11851,
       n_11852;
  wire n_11853, n_11854, n_11855, n_11856, n_11857, n_11858, n_11859,
       n_11860;
  wire n_11861, n_11862, n_11863, n_11864, n_11865, n_11866, n_11867,
       n_11868;
  wire n_11869, n_11870, n_11871, n_11872, n_11873, n_11874, n_11875,
       n_11876;
  wire n_11877, n_11878, n_11879, n_11880, n_11881, n_11882, n_11883,
       n_11884;
  wire n_11885, n_11886, n_11887, n_11888, n_11889, n_11890, n_11891,
       n_11892;
  wire n_11893, n_11894, n_11895, n_11896, n_11897, n_11898, n_11899,
       n_11900;
  wire n_11901, n_11902, n_11903, n_11904, n_11905, n_11906, n_11907,
       n_11908;
  wire n_11909, n_11910, n_11911, n_11912, n_11913, n_11914, n_11915,
       n_11916;
  wire n_11917, n_11918, n_11919, n_11920, n_11921, n_11922, n_11923,
       n_11924;
  wire n_11925, n_11926, n_11927, n_11928, n_11929, n_11930, n_11931,
       n_11932;
  wire n_11933, n_11934, n_11935, n_11936, n_11937, n_11938, n_11939,
       n_11940;
  wire n_11941, n_11942, n_11943, n_11944, n_11945, n_11946, n_11947,
       n_11948;
  wire n_11949, n_11950, n_11951, n_11952, n_11953, n_11954, n_11955,
       n_11956;
  wire n_11958, n_11959, n_11960, n_11961, n_11962, n_11963, n_11964,
       n_11965;
  wire n_11966, n_11967, n_11968, n_11969, n_11970, n_11971, n_11972,
       n_11973;
  wire n_11974, n_11975, n_11976, n_11977, n_11978, n_11979, n_11980,
       n_11981;
  wire n_11982, n_11983, n_11984, n_11985, n_11986, n_11987, n_11988,
       n_11989;
  wire n_11990, n_11991, n_11992, n_11993, n_11994, n_11995, n_11996,
       n_11997;
  wire n_11998, n_11999, n_12000, n_12001, n_12003, n_12004, n_12005,
       n_12006;
  wire n_12007, n_12008, n_12009, n_12010, n_12011, n_12012, n_12013,
       n_12014;
  wire n_12015, n_12016, n_12017, n_12018, n_12019, n_12020, n_12021,
       n_12022;
  wire n_12023, n_12024, n_12025, n_12026, n_12027, n_12028, n_12029,
       n_12030;
  wire n_12031, n_12032, n_12033, n_12034, n_12035, n_12036, n_12037,
       n_12038;
  wire n_12039, n_12040, n_12041, n_12042, n_12043, n_12044, n_12045,
       n_12046;
  wire n_12047, n_12048, n_12049, n_12050, n_12051, n_12052, n_12053,
       n_12054;
  wire n_12055, n_12056, n_12057, n_12058, n_12059, n_12060, n_12061,
       n_12062;
  wire n_12063, n_12064, n_12065, n_12066, n_12067, n_12068, n_12069,
       n_12070;
  wire n_12071, n_12072, n_12073, n_12112, n_12113, n_12114, n_12117,
       n_12118;
  wire n_12120, n_12122, n_12124, n_12126, n_12133, n_12138, n_12147,
       n_12148;
  wire n_12149, n_12152, n_12153, n_12168, n_12172, n_12174, n_12175,
       n_12178;
  wire n_12179, n_12180, n_12181, n_12182, n_12186, n_12189, n_12190,
       n_12191;
  wire n_12192, n_12193, n_12196, n_12197, n_12200, n_12202, n_12204,
       n_12205;
  wire n_12207, n_12210, n_12213, n_12214, n_12215, n_12216, n_12218,
       n_12219;
  wire n_12220, n_12221, n_12223, n_12224, n_12225, n_12227, n_12229,
       n_12231;
  wire n_12233, n_12236, n_12237, n_12238, n_12240, n_12242, n_12243,
       n_12244;
  wire n_12245, n_12252, n_12253, n_12254, n_12255, n_12256, n_12257,
       n_12258;
  wire n_12259, n_12261, n_12262, n_12264, n_12265, n_12266, n_12271,
       n_12272;
  wire n_12278, n_12279, n_12280, n_12281, n_12282, n_12283, n_12284,
       n_12285;
  wire n_12286, n_12287, n_12289, n_12291, n_12293, n_12294, n_12295,
       n_12296;
  wire n_12297, n_12299, n_12300, n_12301, n_12302, n_12303, n_12305,
       n_12306;
  wire n_12308, n_12309, n_12310, n_12311, n_12312, n_12313, n_12314,
       n_12316;
  wire n_12317, n_12318, n_12319, n_12320, n_12321, n_12322, n_12323,
       n_12324;
  wire n_12325, n_12326, n_12327, n_12328, n_12329, n_12330, n_12331,
       n_12332;
  wire n_12333, n_12334, n_12335, n_12336, n_12337, n_12338, n_12339,
       n_12340;
  wire n_12349, n_12350, n_12351, n_12352, n_12353, n_12354, n_12355,
       n_12356;
  wire n_12358, n_12359, n_12360, n_12361, n_12362, n_12363, n_12364,
       n_12365;
  wire n_12366, n_12367, n_12368, n_12369, n_12370, n_12371, n_12372,
       n_12373;
  wire n_12374, n_12375, n_12376, n_12377, n_12378, n_12379, n_12380,
       n_12381;
  wire n_12382, n_12383, n_12384, n_12385, n_12386, n_12387, n_12388,
       n_12389;
  wire n_12390, n_12391, n_12392, n_12393, n_12394, n_12395, n_12396,
       n_12397;
  wire n_12398, n_12399, n_12400, n_12401, n_12402, n_12403, n_12404,
       n_12405;
  wire n_12406, n_12407, n_12408, n_12409, n_12410, n_12417, n_12418,
       n_12419;
  wire n_12440, n_12441, n_12442, n_12443, n_12444, n_12445, n_12448,
       n_12457;
  wire n_12458, n_12459, n_12460, n_12467, n_12468, n_12469, n_12472,
       n_12475;
  wire n_12480, n_12481, n_12484, n_12487, n_12490, n_12493, n_12496,
       n_12499;
  wire n_12507, n_12508, n_12517, n_12518, n_12519, n_12520, n_12525,
       n_12526;
  wire n_12531, n_12532, n_12535, n_12538, n_12547, n_12548, n_12549,
       n_12550;
  wire n_12557, n_12558, n_12559, n_12562, n_12565, n_12568, n_12571,
       n_12574;
  wire n_12581, n_12582, n_12583, n_12590, n_12591, n_12592, n_12599,
       n_12600;
  wire n_12601, n_12604, n_12611, n_12612, n_12613, n_12616, n_12619,
       n_12622;
  wire n_12629, n_12630, n_12631, n_12634, n_12637, n_12640, n_12651,
       n_12652;
  wire n_12653, n_12654, n_12655, n_12660, n_12661, n_12664, n_12671,
       n_12672;
  wire n_12673, n_12680, n_12681, n_12682, n_12685, n_12688, n_12691,
       n_12694;
  wire n_12697, n_12700, n_12703, n_12710, n_12711, n_12712, n_12715,
       n_12718;
  wire n_12725, n_12726, n_12727, n_12730, n_12737, n_12739, n_12742,
       n_12745;
  wire n_12748, n_12751, n_12754, n_12757, n_12762, n_12763, n_12766,
       n_12769;
  wire n_12772, n_12775, n_12778, n_12781, n_12786, n_12787, n_12797,
       n_12798;
  wire n_12799, n_12805, n_12814, n_12817, n_12822, n_12823, n_12831,
       n_12839;
  wire n_12840, n_12841, n_12844, n_12847, n_12850, n_12853, n_12856,
       n_12859;
  wire n_12864, n_12865, n_12868, n_12871, n_12874, n_12881, n_12882,
       n_12883;
  wire n_12888, n_12889, n_12894, n_12895, n_12900, n_12901, n_12906,
       n_12907;
  wire n_12912, n_12913, n_12918, n_12919, n_12924, n_12925, n_12930,
       n_12931;
  wire n_12936, n_12937, n_12942, n_12943, n_12948, n_12949, n_12954,
       n_12955;
  wire n_12960, n_12961, n_12966, n_12967, n_12972, n_12973, n_12978,
       n_12979;
  wire n_12984, n_12985, n_12990, n_12991, n_12996, n_12997, n_13002,
       n_13003;
  wire n_13008, n_13009, n_13014, n_13015, n_13020, n_13021, n_13026,
       n_13027;
  wire n_13034, n_13035, n_13036, n_13039, n_13044, n_13045, n_13050,
       n_13051;
  wire n_13056, n_13057, n_13062, n_13063, n_13068, n_13069, n_13074,
       n_13075;
  wire n_13080, n_13081, n_13086, n_13087, n_13092, n_13093, n_13096,
       n_13099;
  wire n_13104, n_13105, n_13108, n_13111, n_13114, n_13119, n_13120,
       n_13125;
  wire n_13126, n_13131, n_13132, n_13137, n_13138, n_13143, n_13144,
       n_13149;
  wire n_13150, n_13155, n_13156, n_13161, n_13162, n_13167, n_13168,
       n_13173;
  wire n_13174, n_13179, n_13180, n_13185, n_13186, n_13191, n_13192,
       n_13197;
  wire n_13198, n_13203, n_13204, n_13209, n_13210, n_13215, n_13216,
       n_13221;
  wire n_13222, n_13227, n_13228, n_13233, n_13234, n_13239, n_13240,
       n_13245;
  wire n_13246, n_13251, n_13252, n_13257, n_13258, n_13263, n_13264,
       n_13269;
  wire n_13270, n_13275, n_13276, n_13281, n_13282, n_13287, n_13288,
       n_13293;
  wire n_13294, n_13299, n_13300, n_13305, n_13306, n_13311, n_13312,
       n_13317;
  wire n_13318, n_13323, n_13324, n_13329, n_13330, n_13335, n_13336,
       n_13341;
  wire n_13342, n_13347, n_13348, n_13353, n_13354, n_13359, n_13360,
       n_13365;
  wire n_13366, n_13371, n_13372, n_13377, n_13378, n_13383, n_13384,
       n_13389;
  wire n_13390, n_13395, n_13396, n_13401, n_13402, n_13407, n_13408,
       n_13413;
  wire n_13414, n_13419, n_13420, n_13425, n_13426, n_13431, n_13432,
       n_13437;
  wire n_13438, n_13443, n_13444, n_13449, n_13450, n_13483, n_13484,
       n_13485;
  wire n_13486, n_13487, n_13488, n_13489, n_13490, n_13491, n_13492,
       n_13493;
  wire n_13494, n_13495, n_13496, n_13497, n_13498, n_13531, n_13532,
       n_13533;
  wire n_13534, n_13535, n_13536, n_13537, n_13538, n_13539, n_13540,
       n_13541;
  wire n_13542, n_13543, n_13544, n_13545, n_13546, n_13579, n_13580,
       n_13581;
  wire n_13582, n_13583, n_13584, n_13585, n_13586, n_13587, n_13588,
       n_13589;
  wire n_13590, n_13591, n_13592, n_13593, n_13594, n_13627, n_13628,
       n_13629;
  wire n_13630, n_13631, n_13632, n_13633, n_13634, n_13635, n_13636,
       n_13637;
  wire n_13638, n_13639, n_13640, n_13641, n_13642, n_13675, n_13676,
       n_13677;
  wire n_13678, n_13679, n_13680, n_13681, n_13682, n_13683, n_13684,
       n_13685;
  wire n_13686, n_13687, n_13688, n_13689, n_13690, n_13723, n_13724,
       n_13725;
  wire n_13726, n_13727, n_13728, n_13729, n_13730, n_13731, n_13732,
       n_13733;
  wire n_13734, n_13735, n_13736, n_13737, n_13738, n_13771, n_13772,
       n_13773;
  wire n_13774, n_13775, n_13776, n_13777, n_13778, n_13779, n_13780,
       n_13781;
  wire n_13782, n_13783, n_13784, n_13785, n_13786, n_13819, n_13820,
       n_13821;
  wire n_13822, n_13823, n_13824, n_13825, n_13826, n_13827, n_13828,
       n_13829;
  wire n_13830, n_13831, n_13832, n_13833, n_13834, n_13867, n_13868,
       n_13869;
  wire n_13870, n_13871, n_13872, n_13873, n_13874, n_13875, n_13876,
       n_13877;
  wire n_13878, n_13879, n_13880, n_13881, n_13882, n_13915, n_13916,
       n_13917;
  wire n_13918, n_13919, n_13920, n_13921, n_13922, n_13923, n_13924,
       n_13925;
  wire n_13926, n_13927, n_13928, n_13929, n_13930, n_13963, n_13964,
       n_13965;
  wire n_13966, n_13967, n_13968, n_13969, n_13970, n_13971, n_13972,
       n_13973;
  wire n_13974, n_13975, n_13976, n_13977, n_13978, n_14011, n_14012,
       n_14013;
  wire n_14014, n_14015, n_14016, n_14017, n_14018, n_14019, n_14020,
       n_14021;
  wire n_14022, n_14023, n_14024, n_14025, n_14026, n_14059, n_14060,
       n_14061;
  wire n_14062, n_14063, n_14064, n_14065, n_14066, n_14067, n_14068,
       n_14069;
  wire n_14070, n_14071, n_14072, n_14073, n_14074, n_14107, n_14108,
       n_14109;
  wire n_14110, n_14111, n_14112, n_14113, n_14114, n_14115, n_14116,
       n_14117;
  wire n_14118, n_14119, n_14120, n_14121, n_14122, n_14155, n_14156,
       n_14157;
  wire n_14158, n_14159, n_14160, n_14161, n_14162, n_14163, n_14164,
       n_14165;
  wire n_14166, n_14167, n_14168, n_14169, n_14170, n_14203, n_14204,
       n_14205;
  wire n_14206, n_14207, n_14208, n_14209, n_14210, n_14211, n_14212,
       n_14213;
  wire n_14214, n_14215, n_14216, n_14217, n_14218, n_14251, n_14252,
       n_14253;
  wire n_14254, n_14255, n_14256, n_14257, n_14258, n_14259, n_14260,
       n_14261;
  wire n_14262, n_14263, n_14264, n_14265, n_14266, n_14295, n_14296,
       n_14297;
  wire n_14298, n_14299, n_14300, n_14301, n_14302, n_14303, n_14304,
       n_14305;
  wire n_14306, n_14307, n_14308, n_14316, n_14317, n_14322, n_14323,
       n_14328;
  wire n_14329, n_14334, n_14335, n_14340, n_14341, n_14346, n_14347,
       n_14352;
  wire n_14353, n_14358, n_14359, n_14364, n_14365, n_14370, n_14371,
       n_14376;
  wire n_14377, n_14384, n_14385, n_14386, n_14389, n_14394, n_14395,
       n_14402;
  wire n_14404, n_14411, n_14412, n_14413, n_14434, n_14441, n_14442,
       n_14443;
  wire n_14448, n_14449, n_14454, n_14455, n_14458, n_14467, n_14468,
       n_14469;
  wire n_14470, n_14475, n_14476, n_14484, n_14492, n_14493, n_14494,
       n_14508;
  wire n_14509, n_14514, n_14515, n_14520, n_14521, n_14526, n_14527,
       n_14532;
  wire n_14533, n_14538, n_14539, n_14544, n_14545, n_14550, n_14551,
       n_14556;
  wire n_14557, n_14562, n_14563, n_14568, n_14569, n_14574, n_14575,
       n_14583;
  wire n_14584, n_14589, n_14590, n_14595, n_14596, n_14601, n_14602,
       n_14616;
  wire n_14617, n_14625, n_14626, n_14631, n_14632, n_14635, n_14640,
       n_14641;
  wire n_14646, n_14647, n_14652, n_14653, n_14660, n_14661, n_14662,
       n_14667;
  wire n_14668, n_14673, n_14674, n_14679, n_14680, n_14685, n_14686,
       n_14691;
  wire n_14692, n_14697, n_14698, n_14703, n_14704, n_14711, n_14712,
       n_14713;
  wire n_14716, n_14727, n_14728, n_14729, n_14730, n_14731, n_14736,
       n_14737;
  wire n_14742, n_14743, n_14748, n_14749, n_14754, n_14755, n_14760,
       n_14761;
  wire n_14766, n_14767, n_14772, n_14773, n_14778, n_14779, n_14784,
       n_14785;
  wire n_14790, n_14791, n_14796, n_14797, n_14800, n_14803, n_14808,
       n_14809;
  wire n_14816, n_14817, n_14818, n_14825, n_14826, n_14827, n_14830,
       n_14835;
  wire n_14836, n_14841, n_14842, n_14853, n_14854, n_14855, n_14856,
       n_14857;
  wire n_14862, n_14863, n_14868, n_14869, n_14874, n_14875, n_14880,
       n_14881;
  wire n_14886, n_14887, n_14892, n_14893, n_14898, n_14899, n_14904,
       n_14905;
  wire n_14910, n_14911, n_14916, n_14917, n_14920, n_14931, n_14932,
       n_14933;
  wire n_14934, n_14935, n_14940, n_14941, n_14946, n_14947, n_14952,
       n_14953;
  wire n_14958, n_14959, n_14964, n_14965, n_14970, n_14971, n_14976,
       n_14977;
  wire n_14982, n_14983, n_14988, n_14989, n_14992, n_14997, n_14998,
       n_15005;
  wire n_15006, n_15007, n_15012, n_15013, n_15020, n_15021, n_15022,
       n_15025;
  wire n_15030, n_15031, n_15036, n_15037, n_15042, n_15043, n_15046,
       n_15051;
  wire n_15052, n_15055, n_15060, n_15061, n_15066, n_15067, n_15078,
       n_15079;
  wire n_15080, n_15081, n_15082, n_15087, n_15088, n_15093, n_15094,
       n_15099;
  wire n_15100, n_15105, n_15106, n_15111, n_15112, n_15117, n_15118,
       n_15123;
  wire n_15124, n_15129, n_15130, n_15137, n_15138, n_15139, n_15144,
       n_15145;
  wire n_15148, n_15151, n_15154, n_15157, n_15162, n_15163, n_15174,
       n_15175;
  wire n_15176, n_15177, n_15178, n_15183, n_15184, n_15189, n_15190,
       n_15195;
  wire n_15196, n_15201, n_15202, n_15207, n_15208, n_15213, n_15214,
       n_15219;
  wire n_15220, n_15225, n_15226, n_15233, n_15234, n_15235, n_15240,
       n_15241;
  wire n_15244, n_15247, n_15258, n_15259, n_15260, n_15261, n_15262,
       n_15267;
  wire n_15268, n_15273, n_15274, n_15279, n_15280, n_15285, n_15286,
       n_15291;
  wire n_15292, n_15297, n_15298, n_15303, n_15304, n_15309, n_15310,
       n_15317;
  wire n_15318, n_15319, n_15324, n_15325, n_15340, n_15341, n_15342,
       n_15343;
  wire n_15344, n_15345, n_15346, n_15351, n_15352, n_15357, n_15358,
       n_15363;
  wire n_15364, n_15369, n_15370, n_15375, n_15376, n_15381, n_15382,
       n_15387;
  wire n_15388, n_15393, n_15394, n_15397, n_15400, n_15403, n_15406,
       n_15413;
  wire n_15414, n_15415, n_15420, n_15421, n_15426, n_15427, n_15432,
       n_15433;
  wire n_15438, n_15439, n_15444, n_15445, n_15450, n_15451, n_15456,
       n_15457;
  wire n_15462, n_15463, n_15468, n_15469, n_15474, n_15475, n_15480,
       n_15481;
  wire n_15486, n_15487, n_15492, n_15493, n_15498, n_15499, n_15504,
       n_15505;
  wire n_15510, n_15511, n_15514, n_15519, n_15520, n_15525, n_15526,
       n_15531;
  wire n_15532, n_15537, n_15538, n_15543, n_15544, n_15549, n_15550,
       n_15555;
  wire n_15556, n_15561, n_15562, n_15567, n_15568, n_15573, n_15574,
       n_15579;
  wire n_15580, n_15585, n_15586, n_15591, n_15592, n_15597, n_15598,
       n_15603;
  wire n_15604, n_15609, n_15610, n_15615, n_15616, n_15623, n_15624,
       n_15625;
  wire n_15630, n_15631, n_15636, n_15637, n_15642, n_15643, n_15648,
       n_15649;
  wire n_15654, n_15655, n_15660, n_15661, n_15666, n_15667, n_15672,
       n_15673;
  wire n_15678, n_15679, n_15684, n_15685, n_15690, n_15691, n_15696,
       n_15697;
  wire n_15702, n_15703, n_15708, n_15709, n_15714, n_15715, n_15720,
       n_15721;
  wire n_15724, n_15727, n_15730, n_15733, n_15736, n_15739, n_15742,
       n_15745;
  wire n_15748, n_15751, n_15754, n_15757, n_15760, n_15763, n_15766,
       n_15769;
  wire n_15772, n_15775, n_15778, n_15781, n_15784, n_15787, n_15790,
       n_15793;
  wire n_15796, n_15799, n_15802, n_15805, n_15808, n_15811, n_15814,
       n_15817;
  wire n_15820, n_15823, n_15826, n_16180, n_16181, n_16182, n_16183,
       n_16186;
  wire n_16187, n_16188, n_16189, n_16190, n_16191, n_16192, n_16193,
       n_16194;
  wire n_16195, n_16198, n_16199, n_16200, n_16201, n_16202, n_16203,
       n_16204;
  wire n_16205, n_16208, n_16209, n_16210, n_16211, n_16212, n_16213,
       n_16216;
  wire n_16217, n_16218, n_16219, n_16220, n_16221, n_16222, n_16223,
       n_16224;
  wire n_16225, n_16226, n_16227, n_16228, n_16229, n_16230, n_16231,
       n_16232;
  wire n_16233, n_16234, n_16235, n_16236, n_16237, n_16238, n_16239,
       n_16240;
  wire n_16241, n_16242, n_16243, n_16244, n_16245, n_16246, n_16247,
       n_16248;
  wire n_16249, n_16250, n_16251, n_16252, n_16253, n_16256, n_16257,
       n_16258;
  wire n_16259, n_16260, n_16261, n_16262, n_16263, n_16264, n_16265,
       n_16266;
  wire n_16267, n_16268, n_16269, n_16270, n_16271, n_16272, n_16273,
       n_16274;
  wire n_16275, n_16276, n_16277, n_16278, n_16279, n_16280, n_16281,
       n_16282;
  wire n_16283, n_16284, n_16285, n_16286, n_16287, n_16288, n_16289,
       n_16290;
  wire n_16291, n_16292, n_16293, n_16294, n_16295, n_16296, n_16297,
       n_16298;
  wire n_16299, n_16300, n_16301, n_16302, n_16303, n_16304, n_16305,
       n_16306;
  wire n_16307, n_16308, n_16309, n_16310, n_16311, n_16312, n_16313,
       n_16314;
  wire n_16315, n_16316, n_16317, n_16318, n_16319, n_16320, n_16321,
       n_16322;
  wire n_16323, n_16324, n_16325, n_16326, n_16327, n_16328, n_16329,
       n_16330;
  wire n_16331, n_16332, n_16333, n_16334, n_16335, n_16336, n_16337,
       n_16338;
  wire n_16339, n_16340, n_16341, n_16342, n_16343, n_16344, n_16345,
       n_16346;
  wire n_16347, n_16348, n_16349, n_16350, n_16351, n_16352, n_16353,
       n_16354;
  wire n_16355, n_16356, n_16357, n_16358, n_16359, n_16360, n_16361,
       n_16362;
  CDN_flop \data_stack_mem_reg[0][0] (.clk (clk), .d (n_11897), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [0]));
  CDN_flop \data_stack_mem_reg[0][1] (.clk (clk), .d (n_11898), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [1]));
  CDN_flop \data_stack_mem_reg[0][2] (.clk (clk), .d (n_11899), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [2]));
  CDN_flop \data_stack_mem_reg[0][3] (.clk (clk), .d (n_11900), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [3]));
  CDN_flop \data_stack_mem_reg[0][4] (.clk (clk), .d (n_11901), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [4]));
  CDN_flop \data_stack_mem_reg[0][5] (.clk (clk), .d (n_11902), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [5]));
  CDN_flop \data_stack_mem_reg[0][6] (.clk (clk), .d (n_11903), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [6]));
  CDN_flop \data_stack_mem_reg[0][7] (.clk (clk), .d (n_11904), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [7]));
  CDN_flop \data_stack_mem_reg[1][0] (.clk (clk), .d (n_11892), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [0]));
  CDN_flop \data_stack_mem_reg[1][1] (.clk (clk), .d (n_11891), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [1]));
  CDN_flop \data_stack_mem_reg[1][2] (.clk (clk), .d (n_11890), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [2]));
  CDN_flop \data_stack_mem_reg[1][3] (.clk (clk), .d (n_11889), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [3]));
  CDN_flop \data_stack_mem_reg[1][4] (.clk (clk), .d (n_11888), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [4]));
  CDN_flop \data_stack_mem_reg[1][5] (.clk (clk), .d (n_11887), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [5]));
  CDN_flop \data_stack_mem_reg[1][6] (.clk (clk), .d (n_11886), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [6]));
  CDN_flop \data_stack_mem_reg[1][7] (.clk (clk), .d (n_11885), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [7]));
  CDN_flop \data_stack_mem_reg[2][0] (.clk (clk), .d (n_11920), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [0]));
  CDN_flop \data_stack_mem_reg[2][1] (.clk (clk), .d (n_11914), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [1]));
  CDN_flop \data_stack_mem_reg[2][2] (.clk (clk), .d (n_11915), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [2]));
  CDN_flop \data_stack_mem_reg[2][3] (.clk (clk), .d (n_11916), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [3]));
  CDN_flop \data_stack_mem_reg[2][4] (.clk (clk), .d (n_11918), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [4]));
  CDN_flop \data_stack_mem_reg[2][5] (.clk (clk), .d (n_11917), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [5]));
  CDN_flop \data_stack_mem_reg[2][6] (.clk (clk), .d (n_11919), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [6]));
  CDN_flop \data_stack_mem_reg[2][7] (.clk (clk), .d (n_11921), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [7]));
  CDN_flop \data_stack_mem_reg[3][0] (.clk (clk), .d (n_11875), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [0]));
  CDN_flop \data_stack_mem_reg[3][1] (.clk (clk), .d (n_11877), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [1]));
  CDN_flop \data_stack_mem_reg[3][2] (.clk (clk), .d (n_11878), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [2]));
  CDN_flop \data_stack_mem_reg[3][3] (.clk (clk), .d (n_11879), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [3]));
  CDN_flop \data_stack_mem_reg[3][4] (.clk (clk), .d (n_11874), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [4]));
  CDN_flop \data_stack_mem_reg[3][5] (.clk (clk), .d (n_11876), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [5]));
  CDN_flop \data_stack_mem_reg[3][6] (.clk (clk), .d (n_11880), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [6]));
  CDN_flop \data_stack_mem_reg[3][7] (.clk (clk), .d (n_11873), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [7]));
  CDN_flop \data_stack_mem_reg[4][0] (.clk (clk), .d (n_12052), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [0]));
  CDN_flop \data_stack_mem_reg[4][1] (.clk (clk), .d (n_12051), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [1]));
  CDN_flop \data_stack_mem_reg[4][2] (.clk (clk), .d (n_12050), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [2]));
  CDN_flop \data_stack_mem_reg[4][3] (.clk (clk), .d (n_12048), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [3]));
  CDN_flop \data_stack_mem_reg[4][4] (.clk (clk), .d (n_12049), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [4]));
  CDN_flop \data_stack_mem_reg[4][5] (.clk (clk), .d (n_12046), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [5]));
  CDN_flop \data_stack_mem_reg[4][6] (.clk (clk), .d (n_12047), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [6]));
  CDN_flop \data_stack_mem_reg[4][7] (.clk (clk), .d (n_12045), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [7]));
  CDN_flop \data_stack_mem_reg[5][0] (.clk (clk), .d (n_11978), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [0]));
  CDN_flop \data_stack_mem_reg[5][1] (.clk (clk), .d (n_11972), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [1]));
  CDN_flop \data_stack_mem_reg[5][2] (.clk (clk), .d (n_11977), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [2]));
  CDN_flop \data_stack_mem_reg[5][3] (.clk (clk), .d (n_11979), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [3]));
  CDN_flop \data_stack_mem_reg[5][4] (.clk (clk), .d (n_11974), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [4]));
  CDN_flop \data_stack_mem_reg[5][5] (.clk (clk), .d (n_11976), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [5]));
  CDN_flop \data_stack_mem_reg[5][6] (.clk (clk), .d (n_11975), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [6]));
  CDN_flop \data_stack_mem_reg[5][7] (.clk (clk), .d (n_11973), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [7]));
  CDN_flop \data_stack_mem_reg[6][0] (.clk (clk), .d (n_11983), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [0]));
  CDN_flop \data_stack_mem_reg[6][1] (.clk (clk), .d (n_11987), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [1]));
  CDN_flop \data_stack_mem_reg[6][2] (.clk (clk), .d (n_11988), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [2]));
  CDN_flop \data_stack_mem_reg[6][3] (.clk (clk), .d (n_11989), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [3]));
  CDN_flop \data_stack_mem_reg[6][4] (.clk (clk), .d (n_11984), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [4]));
  CDN_flop \data_stack_mem_reg[6][5] (.clk (clk), .d (n_11985), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [5]));
  CDN_flop \data_stack_mem_reg[6][6] (.clk (clk), .d (n_11986), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [6]));
  CDN_flop \data_stack_mem_reg[6][7] (.clk (clk), .d (n_11990), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [7]));
  CDN_flop \data_stack_mem_reg[7][0] (.clk (clk), .d (n_11997), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [0]));
  CDN_flop \data_stack_mem_reg[7][1] (.clk (clk), .d (n_11994), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [1]));
  CDN_flop \data_stack_mem_reg[7][2] (.clk (clk), .d (n_12000), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [2]));
  CDN_flop \data_stack_mem_reg[7][3] (.clk (clk), .d (n_11999), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [3]));
  CDN_flop \data_stack_mem_reg[7][4] (.clk (clk), .d (n_11998), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [4]));
  CDN_flop \data_stack_mem_reg[7][5] (.clk (clk), .d (n_11995), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [5]));
  CDN_flop \data_stack_mem_reg[7][6] (.clk (clk), .d (n_11996), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [6]));
  CDN_flop \data_stack_mem_reg[7][7] (.clk (clk), .d (n_11993), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [7]));
  CDN_flop \data_stack_mem_reg[8][0] (.clk (clk), .d (n_11491), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [0]));
  CDN_flop \data_stack_mem_reg[8][1] (.clk (clk), .d (n_11487), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [1]));
  CDN_flop \data_stack_mem_reg[8][2] (.clk (clk), .d (n_11492), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [2]));
  CDN_flop \data_stack_mem_reg[8][3] (.clk (clk), .d (n_11488), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [3]));
  CDN_flop \data_stack_mem_reg[8][4] (.clk (clk), .d (n_11494), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [4]));
  CDN_flop \data_stack_mem_reg[8][5] (.clk (clk), .d (n_11489), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [5]));
  CDN_flop \data_stack_mem_reg[8][6] (.clk (clk), .d (n_11493), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [6]));
  CDN_flop \data_stack_mem_reg[8][7] (.clk (clk), .d (n_11490), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [7]));
  CDN_flop \data_stack_pointer_reg[0] (.clk (clk), .d (n_12026), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[0]));
  CDN_flop \data_stack_pointer_reg[1] (.clk (clk), .d (n_12025), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[1]));
  CDN_flop \data_stack_pointer_reg[2] (.clk (clk), .d (n_11952), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[2]));
  CDN_flop \data_stack_pointer_reg[3] (.clk (clk), .d (n_12027), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[3]));
  CDN_flop dout_valid_reg(.clk (clk), .d (n_11479), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (dout_valid));
  or g14025 (n_11532, out_fifo_write_pointer[1],
       out_fifo_write_pointer[0]);
  nand g18391 (n_11512, data_stack_pointer[1], data_stack_pointer[0]);
  nand g18413 (n_11518, \data_stack_mem[1] [0], \data_stack_mem[0] [0]);
  nand g18426 (n_11566, n_11528, \data_stack_mem[7] [0]);
  nand g18430 (n_11573, n_11524, \data_stack_mem[3] [0]);
  nand g18434 (n_11571, n_11525, \data_stack_mem[4] [0]);
  nand g18438 (n_11569, n_11526, \data_stack_mem[5] [0]);
  nand g18442 (n_11574, n_11523, \data_stack_mem[2] [0]);
  nand g18446 (n_11568, n_11527, \data_stack_mem[6] [0]);
  or g18455 (n_11483, data_stack_pointer[2], n_11482);
  or g18712 (n_11475, sh_bit_cnt[0], sh_bit_cnt[1]);
  nand g18750 (n_11565, n_11529, \data_stack_mem[8] [0]);
  or g18774 (n_11455, n_11454, sh_reg_out_bit_counter[3]);
  or g18775 (n_11456, n_11455, sh_reg_out_bit_counter[4]);
  or g18778 (n_11503, data_stack_pointer[2], data_stack_pointer[1]);
  or g18786 (n_11453, sh_reg_out_bit_counter[0],
       sh_reg_out_bit_counter[1]);
  or g18787 (n_11454, n_11453, sh_reg_out_bit_counter[2]);
  or g18802 (n_11514, data_stack_pointer[3], data_stack_pointer[1]);
  or g18809 (n_11555, n_11532, n_11497);
  not g18811 (n_11941, n_11555);
  or g18815 (n_11547, n_11546, n_11533);
  not g18817 (n_11942, n_11547);
  or g18819 (n_11551, n_11538, n_11533);
  not g18821 (n_11943, n_11551);
  or g18823 (n_11559, n_11546, n_11497);
  not g18825 (n_11944, n_11559);
  or g18827 (n_11534, n_11532, n_11533);
  not g18829 (n_11945, n_11534);
  or g18831 (n_11539, n_11538, n_11497);
  not g18833 (n_11946, n_11539);
  or g19130 (n_11968, data_stack_pointer[3], wc);
  not gc (wc, data_stack_pointer[2]);
  not g22670 (n_11462, rst_n);
  not g22671 (n_11463, enable_n);
  or g22688 (n_11509, n_11508, data_stack_pointer[0]);
  or g22692 (n_11538, wc0, out_fifo_write_pointer[0]);
  not gc0 (wc0, out_fifo_write_pointer[1]);
  or g22693 (n_11546, out_fifo_write_pointer[1], wc1);
  not gc1 (wc1, out_fifo_write_pointer[0]);
  nand g22726 (n_12001, out_fifo_read_pointer[1],
       out_fifo_read_pointer[0]);
  or g22903 (n_11481, n_11476, sh_bit_cnt[3]);
  or g22953 (n_11905, n_11481, wc2);
  not gc2 (wc2, sh_reg_in[8]);
  or g23102 (n_11533, n_11905, out_fifo_write_pointer[2]);
  or g23170 (n_11497, n_11905, wc3);
  not gc3 (wc3, out_fifo_write_pointer[2]);
  or g23297 (n_12147, n_11516, \data_stack_mem[4] [2]);
  or g23369 (n_12178, n_11742, \data_stack_mem[2] [6]);
  or g23372 (n_12179, n_11704, \data_stack_mem[3] [5]);
  or g23375 (n_12180, n_11677, \data_stack_mem[3] [4]);
  nand g23378 (n_12181, n_11764, \data_stack_mem[3] [7]);
  or g23381 (n_12182, n_11601, \data_stack_mem[5] [2]);
  or g23398 (n_12189, n_11599, \data_stack_mem[6] [2]);
  or g23401 (n_12190, n_11611, \data_stack_mem[4] [2]);
  nand g23407 (n_12192, data_stack_pointer[3], \data_stack_mem[7] [0]);
  or g23410 (n_12193, n_11734, \data_stack_mem[7] [6]);
  or g23418 (n_12196, n_11672, \data_stack_mem[2] [4]);
  nand g23441 (n_12205, n_11759, \data_stack_mem[7] [7]);
  or g23446 (n_12207, n_11698, \data_stack_mem[7] [5]);
  or g23460 (n_12213, n_11606, \data_stack_mem[1] [2]);
  or g23463 (n_12214, n_11706, \data_stack_mem[2] [5]);
  or g23466 (n_12215, n_11643, \data_stack_mem[1] [3]);
  or g23469 (n_12216, n_11642, \data_stack_mem[2] [3]);
  or g23481 (n_12220, n_11635, \data_stack_mem[6] [3]);
  or g23484 (n_12221, n_11637, \data_stack_mem[5] [3]);
  or g23492 (n_12224, n_11597, \data_stack_mem[7] [2]);
  or g23506 (n_12229, n_11702, \data_stack_mem[4] [5]);
  or g23527 (n_12237, n_11665, \data_stack_mem[7] [4]);
  or g23535 (n_12240, n_11700, \data_stack_mem[6] [5]);
  nand g23543 (n_12243, n_11774, \data_stack_mem[6] [7]);
  or g23546 (n_12244, n_11604, \data_stack_mem[2] [2]);
  or g23569 (n_12253, n_11481, sh_reg_in[8]);
  or g23570 (n_11482, n_12253, data_stack_pointer[1]);
  nand g23575 (n_12255, n_11766, \data_stack_mem[2] [7]);
  or g23577 (n_11767, wc4, n_12218);
  not gc4 (wc4, n_12255);
  or g23578 (n_12256, n_11633, \data_stack_mem[7] [3]);
  or g23581 (n_12257, n_11582, \data_stack_mem[8] [1]);
  nand g23600 (n_12264, n_11760, \data_stack_mem[5] [7]);
  or g23602 (n_11761, wc5, n_12227);
  not gc5 (wc5, n_12264);
  nand g23603 (n_12265, n_11762, \data_stack_mem[4] [7]);
  or g23605 (n_11763, wc6, n_12258);
  not gc6 (wc6, n_12265);
  nand g23606 (n_12266, n_11517, \data_stack_mem[2] [0]);
  or g23619 (n_12271, n_11738, \data_stack_mem[4] [6]);
  or g23622 (n_12272, n_11740, \data_stack_mem[3] [6]);
  or g23646 (n_12191, wc7, \data_stack_mem[1] [1]);
  not gc7 (wc7, n_11518);
  or g23647 (n_12262, n_11516, wc8);
  not gc8 (wc8, \data_stack_mem[4] [0]);
  or g23662 (n_12133, wc9, \data_stack_mem[2] [3]);
  not gc9 (wc9, n_11517);
  or g23704 (n_12238, wc10, \data_stack_mem[4] [1]);
  not gc10 (wc10, n_11571);
  or g23710 (n_12225, wc11, \data_stack_mem[5] [1]);
  not gc11 (wc11, n_11569);
  or g23727 (n_12259, wc12, \data_stack_mem[7] [1]);
  not gc12 (wc12, n_11566);
  or g23785 (n_11765, n_12223, wc13);
  not gc13 (wc13, n_12181);
  or g23811 (n_11817, wc14, n_11777);
  not gc14 (wc14, n_11788);
  or g23829 (n_11790, wc15, n_12202);
  not gc15 (wc15, n_12205);
  or g23999 (n_12278, \data_stack_mem[3] [1], wc16);
  not gc16 (wc16, n_11573);
  nand g24001 (n_12279, \data_stack_mem[1] [0], n_11508);
  or g24007 (n_12281, \data_stack_mem[8] [7], n_11791);
  or g24009 (n_12282, \data_stack_mem[6] [4], n_11680);
  or g24011 (n_12283, \data_stack_mem[4] [3], n_11639);
  or g24013 (n_12284, \data_stack_mem[5] [4], n_11679);
  or g24018 (n_12286, \data_stack_mem[5] [5], n_11712);
  or g24032 (n_12293, \data_stack_mem[3] [3], n_11641);
  or g24034 (n_12294, \data_stack_mem[6] [6], n_11750);
  or g24036 (n_12295, wc17, \data_stack_mem[2] [1]);
  not gc17 (wc17, n_11574);
  or g24038 (n_12296, \data_stack_mem[4] [4], n_11670);
  or g24040 (n_12297, \data_stack_mem[3] [2], n_11602);
  or g24048 (n_12301, \data_stack_mem[8] [6], n_11732);
  or g24050 (n_12302, \data_stack_mem[8] [7], n_11504);
  or g24062 (n_12308, \data_stack_mem[8] [5], n_11716);
  or g24066 (n_12310, \data_stack_mem[8] [6], n_11504);
  or g24070 (n_12312, \data_stack_mem[5] [6], n_11748);
  or g24078 (n_12316, wc18, \data_stack_mem[6] [1]);
  not gc18 (wc18, n_11568);
  or g24080 (n_12317, \data_stack_mem[8] [4], n_11684);
  or g24084 (n_12319, \data_stack_mem[8] [5], n_11504);
  or g24088 (n_12321, \data_stack_mem[8] [3], n_11631);
  or g24090 (n_12322, \data_stack_mem[8] [2], n_11617);
  or g24092 (n_12323, \data_stack_mem[0] [4], \data_stack_mem[1] [4]);
  or g24096 (n_12325, \data_stack_mem[8] [4], n_11504);
  or g24100 (n_12327, \data_stack_mem[0] [5], \data_stack_mem[1] [5]);
  or g24102 (n_12328, \data_stack_mem[0] [6], \data_stack_mem[1] [6]);
  or g24106 (n_12330, wc19, data_stack_pointer[3]);
  not gc19 (wc19, n_11512);
  or g24108 (n_12331, wc20, data_stack_pointer[2]);
  not gc20 (wc20, data_stack_pointer[0]);
  or g24116 (n_12335, \data_stack_mem[8] [2], n_11504);
  or g24124 (n_12339, \data_stack_mem[8] [3], n_11504);
  or g24146 (n_12350, \data_stack_mem[8] [1], n_11504);
  or g24150 (n_12352, \data_stack_mem[0] [7], \data_stack_mem[1] [7]);
  or g24170 (n_12362, n_11469, n_12001);
  nand g24180 (n_12367, data_stack_pointer[3], n_11503);
  or g24188 (n_12371, \data_stack_mem[2] [0], wc21);
  not gc21 (wc21, n_11517);
  or g24192 (n_12373, \data_stack_mem[4] [0], n_11516);
  or g24196 (n_12375, \data_stack_mem[8] [0], n_11504);
  or g24204 (n_12379, \data_stack_mem[4] [6], n_11516);
  or g24208 (n_12381, \data_stack_mem[2] [6], wc22);
  not gc22 (wc22, n_11517);
  or g24210 (n_12382, \data_stack_mem[4] [1], n_11516);
  or g24212 (n_12383, \data_stack_mem[1] [1], wc23);
  not gc23 (wc23, n_11508);
  or g24214 (n_12384, \data_stack_mem[2] [1], wc24);
  not gc24 (wc24, n_11517);
  or g24220 (n_12387, \data_stack_mem[4] [4], n_11516);
  or g24224 (n_12389, \data_stack_mem[2] [5], wc25);
  not gc25 (wc25, n_11517);
  or g24228 (n_12391, \data_stack_mem[2] [4], wc26);
  not gc26 (wc26, n_11517);
  or g24232 (n_12393, \data_stack_mem[4] [5], n_11516);
  or g24244 (n_12399, \data_stack_mem[4] [7], n_11516);
  or g24248 (n_12401, \data_stack_mem[2] [7], wc27);
  not gc27 (wc27, n_11517);
  or g24250 (n_12402, \data_stack_mem[1] [2], wc28);
  not gc28 (wc28, n_11508);
  or g24252 (n_12403, \data_stack_mem[2] [2], wc29);
  not gc29 (wc29, n_11517);
  or g24262 (n_12408, \data_stack_mem[1] [3], wc30);
  not gc30 (wc30, n_11508);
  or g24264 (n_12409, \data_stack_mem[4] [3], n_11516);
  or g24285 (n_12329, n_12440, n_12441);
  nand g26500 (n_12020, n_15702, n_15703);
  nand g26501 (n_12019, n_15696, n_15697);
  nand g26502 (n_12015, n_15678, n_15679);
  nand g26503 (n_12022, n_15714, n_15715);
  nand g26504 (n_12018, n_15720, n_15721);
  nand g26505 (n_12021, n_15708, n_15709);
  nand g26506 (n_12016, n_15684, n_15685);
  nand g26507 (n_12017, n_15690, n_15691);
  or g26511 (n_15721, wc31, n_11544);
  not gc31 (wc31, n_12014);
  or g26515 (n_15679, wc32, n_11500);
  not gc32 (wc32, n_12014);
  nand g26516 (n_11929, n_15630, n_15631);
  nand g26517 (n_11853, n_15567, n_15568);
  nand g26518 (n_11938, n_15654, n_15655);
  nand g26519 (n_11857, n_15585, n_15586);
  nand g26520 (n_11856, n_15615, n_15616);
  nand g26521 (n_11936, n_15648, n_15649);
  nand g26522 (n_11859, n_15597, n_15598);
  or g26523 (n_16180, wc33, n_11925);
  not gc33 (wc33, n_12013);
  or g26524 (n_16181, n_12013, wc34);
  not gc34 (wc34, n_11925);
  nand g26525 (n_12014, n_16180, n_16181);
  nand g26526 (n_11934, n_15642, n_15643);
  nand g26527 (n_11854, n_15573, n_15574);
  nand g26528 (n_11932, n_15672, n_15673);
  nand g26529 (n_11858, n_15591, n_15592);
  nand g26530 (n_11931, n_15636, n_15637);
  nand g26531 (n_11926, n_15666, n_15667);
  nand g26532 (n_11855, n_15579, n_15580);
  nand g26533 (n_11860, n_15603, n_15604);
  nand g26534 (n_11940, n_15660, n_15661);
  nand g26535 (n_11833, n_15525, n_15526);
  nand g26536 (n_11835, n_15531, n_15532);
  nand g26537 (n_11839, n_15537, n_15538);
  nand g26538 (n_11841, n_15543, n_15544);
  nand g26539 (n_11843, n_15549, n_15550);
  nand g26540 (n_11845, n_15555, n_15556);
  nand g26541 (n_11831, n_15561, n_15562);
  or g26542 (n_15568, wc35, n_11500);
  not gc35 (wc35, n_11852);
  nand g26545 (n_12013, n_16182, n_16183);
  nand g26554 (n_11837, n_15609, n_15610);
  or g26555 (n_15616, wc36, n_11544);
  not gc36 (wc36, n_11852);
  nand g26562 (n_11933, n_15468, n_15469);
  nand g26563 (n_11803, n_15432, n_15433);
  nand g26564 (n_11799, n_15426, n_15427);
  nand g26566 (n_11937, n_15480, n_15481);
  nand g26567 (n_11805, n_15438, n_15439);
  nand g26568 (n_11797, n_15420, n_15421);
  or g26569 (n_15610, wc37, n_11544);
  not gc37 (wc37, n_11830);
  nand g26571 (n_11807, n_15444, n_15445);
  nand g26572 (n_11801, n_15510, n_15511);
  nand g26573 (n_11939, n_15486, n_15487);
  nand g26578 (n_11809, n_15450, n_15451);
  nand g26579 (n_11935, n_15474, n_15475);
  nand g26580 (n_12011, n_15498, n_15499);
  nand g26582 (n_11928, n_15456, n_15457);
  nand g26583 (n_11795, n_15504, n_15505);
  nand g26584 (n_11925, n_15624, n_15625);
  nand g26586 (n_11930, n_15462, n_15463);
  or g26587 (n_16186, wc38, n_11851);
  not gc38 (wc38, n_11848);
  or g26588 (n_16187, n_11848, wc39);
  not gc39 (wc39, n_11851);
  nand g26589 (n_11852, n_16186, n_16187);
  or g26590 (n_15562, wc40, n_11500);
  not gc40 (wc40, n_11830);
  nand g26591 (n_12010, n_15492, n_15493);
  nand g26598 (n_11830, n_15519, n_15520);
  nand g26600 (n_11836, n_15393, n_15394);
  or g26601 (n_15457, n_11536, n_11927);
  nand g26602 (n_11816, n_15387, n_15388);
  nand g26603 (n_11844, n_15381, n_15382);
  or g26604 (n_15463, n_11541, n_11927);
  nand g26605 (n_11842, n_15375, n_15376);
  nand g26606 (n_11840, n_15369, n_15370);
  or g26607 (n_15469, n_11549, n_11927);
  nand g26608 (n_11838, n_15363, n_15364);
  nand g26609 (n_11834, n_15357, n_15358);
  or g26610 (n_15475, n_11553, n_11927);
  nand g26611 (n_11832, n_15351, n_15352);
  nand g26612 (n_15625, n_12313, n_11924);
  or g26613 (n_15481, n_11557, n_11927);
  nand g26614 (n_16188, n_11846, n_11847);
  or g26615 (n_16189, n_11846, n_11847);
  nand g26616 (n_11848, n_16188, n_16189);
  or g26618 (n_15486, n_11561, n_11927);
  or g26620 (n_15499, n_11927, n_11544);
  or g26621 (n_15493, n_11927, n_11500);
  or g26623 (n_15352, n_11536, wc41);
  not gc41 (wc41, n_11815);
  or g26624 (n_15364, n_11549, wc42);
  not gc42 (wc42, n_11815);
  or g26625 (n_12313, n_11829, wc43);
  not gc43 (wc43, n_15514);
  or g26626 (n_15381, n_11561, wc44);
  not gc44 (wc44, n_11815);
  or g26627 (n_15624, n_15623, wc45);
  not gc45 (wc45, n_11827);
  or g26628 (n_15358, n_11541, wc46);
  not gc46 (wc46, n_11815);
  or g26629 (n_15376, n_11557, wc47);
  not gc47 (wc47, n_11815);
  nand g26630 (n_11794, n_15414, n_15415);
  nand g26631 (n_15520, n_11827, n_11829);
  or g26632 (n_15394, n_11544, wc48);
  not gc48 (wc48, n_11815);
  or g26633 (n_15370, n_11553, wc49);
  not gc49 (wc49, n_11815);
  nand g26636 (n_11847, n_16190, n_16191);
  or g26637 (n_15388, n_11500, wc50);
  not gc50 (wc50, n_11815);
  or g26640 (n_15623, n_11924, n_11828);
  nand g26641 (n_15415, n_11789, n_12174);
  or g26642 (n_11829, n_12174, wc51);
  not gc51 (wc51, n_15403);
  or g26643 (n_15519, n_11827, n_11828);
  nand g26644 (n_15346, n_15343, n_15344);
  or g26645 (n_15414, n_15413, n_11506);
  or g26646 (n_16192, wc52, n_11656);
  not gc52 (wc52, n_11850);
  or g26647 (n_16193, n_11850, wc53);
  not gc53 (wc53, n_11656);
  nand g26648 (n_11851, n_16192, n_16193);
  nand g26649 (n_12174, n_15397, n_11505);
  or g26650 (n_11828, n_15400, n_11506);
  or g26652 (n_15514, n_11827, n_11502);
  or g26653 (n_16194, wc54, n_11723);
  not gc54 (wc54, n_11849);
  or g26654 (n_16195, n_11849, wc55);
  not gc55 (wc55, n_11723);
  nand g26655 (n_11850, n_16194, n_16195);
  nand g26656 (n_11758, n_15303, n_15304);
  nand g26657 (n_11800, n_15309, n_15310);
  nand g26658 (n_15344, n_11509, n_11811);
  or g26662 (n_15397, n_11502, n_11793);
  nand g26663 (n_11804, n_15285, n_15286);
  nand g26664 (n_11798, n_15273, n_15274);
  nand g26665 (n_11796, n_15267, n_15268);
  nand g26666 (n_11808, n_15297, n_15298);
  nand g26667 (n_11802, n_15279, n_15280);
  nand g26668 (n_15400, n_11793, n_11789);
  nand g26669 (n_11806, n_15291, n_15292);
  or g26670 (n_15280, n_11549, wc56);
  not gc56 (wc56, n_11757);
  or g26671 (n_15268, n_11536, wc57);
  not gc57 (wc57, n_11757);
  or g26672 (n_15310, n_11544, wc58);
  not gc58 (wc58, n_11757);
  or g26673 (n_15304, n_11500, wc59);
  not gc59 (wc59, n_11757);
  nand g26674 (n_16198, n_11817, n_11826);
  or g26675 (n_16199, n_11817, n_11826);
  nand g26676 (n_11827, n_16198, n_16199);
  or g26677 (n_15297, n_11561, wc60);
  not gc60 (wc60, n_11757);
  or g26678 (n_15403, n_11789, n_11502);
  or g26679 (n_15292, n_11557, wc61);
  not gc61 (wc61, n_11757);
  or g26680 (n_15286, n_11553, wc62);
  not gc62 (wc62, n_11757);
  nand g26681 (n_11811, n_15318, n_15319);
  nand g26682 (n_11793, n_15324, n_15325);
  nand g26685 (n_11849, n_16200, n_16201);
  or g26686 (n_15274, n_11541, wc63);
  not gc63 (wc63, n_11757);
  nand g26687 (n_15324, n_12281, n_11792);
  or g26688 (n_15318, n_15317, n_11506);
  nand g26689 (n_16202, n_11777, n_11788);
  or g26690 (n_16203, n_11777, n_11788);
  nand g26691 (n_11789, n_16202, n_16203);
  nand g26693 (n_15262, n_15259, n_15260);
  nand g26695 (n_15319, n_12300, n_11791);
  or g26696 (n_15317, n_11791, wc64);
  not gc64 (wc64, n_11810);
  nand g26697 (n_15325, \data_stack_mem[8] [7], n_11791);
  nand g26698 (n_11725, n_15183, n_15184);
  nand g26699 (n_11727, n_15225, n_15226);
  nand g26700 (n_15260, n_11509, n_11753);
  or g26701 (n_15247, wc65, n_11776);
  not gc65 (wc65, n_12205);
  nand g26702 (n_12300, n_11505, n_15244);
  nand g26703 (n_11724, n_15219, n_15220);
  nand g26704 (n_11731, n_15213, n_15214);
  nand g26705 (n_16204, n_11790, n_11776);
  or g26706 (n_16205, n_11790, n_11776);
  nand g26707 (n_11791, n_16204, n_16205);
  nand g26708 (n_11730, n_15207, n_15208);
  nand g26712 (n_11729, n_15201, n_15202);
  nand g26713 (n_11728, n_15195, n_15196);
  nand g26714 (n_11726, n_15189, n_15190);
  or g26715 (n_15190, n_11541, wc66);
  not gc66 (wc66, n_11723);
  or g26716 (n_15196, n_11549, wc67);
  not gc67 (wc67, n_11723);
  or g26717 (n_15220, n_11500, wc68);
  not gc68 (wc68, n_11723);
  or g26718 (n_15244, n_11506, n_11810);
  nand g26719 (n_16208, n_11818, n_11825);
  or g26720 (n_16209, n_11818, n_11825);
  nand g26721 (n_11826, n_16208, n_16209);
  or g26722 (n_15184, n_11536, wc69);
  not gc69 (wc69, n_11723);
  nand g26723 (n_11753, n_15234, n_15235);
  or g26724 (n_15213, n_11561, wc70);
  not gc70 (wc70, n_11723);
  or g26725 (n_15202, n_11553, wc71);
  not gc71 (wc71, n_11723);
  or g26726 (n_15208, n_11557, wc72);
  not gc72 (wc72, n_11723);
  nand g26727 (n_11776, n_15240, n_15241);
  or g26728 (n_15226, n_11544, wc73);
  not gc73 (wc73, n_11723);
  nand g26732 (n_11810, n_16210, n_16211);
  nand g26734 (n_15235, n_12309, n_11752);
  nand g26735 (n_16212, n_11778, n_11787);
  or g26736 (n_16213, n_11778, n_11787);
  nand g26737 (n_11788, n_16212, n_16213);
  nand g26739 (n_12202, data_stack_pointer[3], n_15151);
  nand g26740 (n_12291, n_15138, n_15139);
  nand g26741 (n_12309, n_11505, n_15154);
  nand g26742 (n_11792, n_15162, n_15163);
  or g26743 (n_11778, n_11775, wc74);
  not gc74 (wc74, n_15157);
  nand g26744 (n_15178, n_15175, n_15176);
  or g26745 (n_15234, n_15233, n_11506);
  nand g26746 (n_15162, n_12301, n_11752);
  nand g26747 (n_11695, n_15105, n_15106);
  or g26749 (n_15154, n_11506, n_11733);
  or g26751 (n_15138, n_15137, n_11513);
  nand g26752 (n_11693, n_15129, n_15130);
  nand g26753 (n_15176, n_11509, n_11719);
  nand g26754 (n_11690, n_15123, n_15124);
  or g26755 (n_15151, \data_stack_mem[7] [7], n_11759);
  nand g26758 (n_11922, n_12168, n_12233);
  nand g26759 (n_11697, n_15117, n_15118);
  nand g26760 (n_11691, n_15087, n_15088);
  nand g26761 (n_11694, n_15099, n_15100);
  nand g26762 (n_11696, n_15111, n_15112);
  nand g26763 (n_11692, n_15093, n_15094);
  or g26764 (n_11775, wc75, n_11513);
  not gc75 (wc75, n_15148);
  nand g26765 (n_16216, n_11735, n_11751);
  or g26766 (n_16217, n_11735, n_11751);
  nand g26767 (n_11752, n_16216, n_16217);
  or g26768 (n_15106, n_11553, wc76);
  not gc76 (wc76, n_11689);
  or g26769 (n_15100, n_11549, wc77);
  not gc77 (wc77, n_11689);
  nand g26772 (n_11733, n_16218, n_16219);
  or g26773 (n_15137, wc78, n_11774);
  not gc78 (wc78, \data_stack_mem[6] [7]);
  or g26774 (n_15094, n_11541, wc79);
  not gc79 (wc79, n_11689);
  or g26775 (n_15112, n_11557, wc80);
  not gc80 (wc80, n_11689);
  or g26776 (n_15117, n_11561, wc81);
  not gc81 (wc81, n_11689);
  or g26777 (n_15088, n_11536, wc82);
  not gc82 (wc82, n_11689);
  or g26778 (n_15130, n_11544, wc83);
  not gc83 (wc83, n_11689);
  nand g26779 (n_11759, n_15051, n_15826);
  nand g26781 (n_16220, n_11819, n_11824);
  or g26782 (n_16221, n_11819, n_11824);
  nand g26783 (n_11825, n_16220, n_16221);
  or g26784 (n_15124, n_11500, wc84);
  not gc84 (wc84, n_11689);
  nand g26785 (n_11719, n_15144, n_15145);
  or g26786 (n_15148, \data_stack_mem[6] [7], n_11774);
  nand g26787 (n_15163, \data_stack_mem[8] [6], n_11732);
  nand g26788 (n_16222, n_11689, n_11622);
  or g26789 (n_16223, n_11689, n_11622);
  nand g26790 (n_11846, n_16222, n_16223);
  nand g26791 (n_15826, n_11751, n_12193);
  or g26792 (n_15144, wc85, n_11506);
  not gc85 (wc85, n_12318);
  nand g26793 (n_11774, n_15060, n_15061);
  nand g26795 (n_16224, n_11779, n_11786);
  or g26796 (n_16225, n_11779, n_11786);
  nand g26797 (n_11787, n_16224, n_16225);
  nand g26798 (n_11732, n_15066, n_15067);
  nand g26799 (n_16226, n_11761, n_11772);
  or g26800 (n_16227, n_11761, n_11772);
  nand g26801 (n_11773, n_16226, n_16227);
  nand g26803 (n_15066, n_12308, n_11718);
  nand g26804 (n_16228, n_11737, n_11750);
  or g26805 (n_16229, n_11737, n_11750);
  nand g26806 (n_11751, n_16228, n_16229);
  or g26807 (n_11779, n_12227, wc86);
  not gc86 (wc86, n_15055);
  nand g26808 (n_15060, n_12294, n_11736);
  nand g26809 (n_15082, n_15079, n_15080);
  or g26810 (n_16230, wc87, n_11718);
  not gc87 (wc87, n_11717);
  or g26811 (n_16231, n_11717, wc88);
  not gc88 (wc88, n_11718);
  nand g26812 (n_12318, n_16230, n_16231);
  nand g26813 (n_15052, n_12193, n_15051);
  nand g26814 (n_15061, \data_stack_mem[6] [6], n_11750);
  or g26815 (n_11737, n_15007, n_11513);
  nand g26818 (n_15051, \data_stack_mem[7] [6], n_11734);
  nand g26820 (n_15080, n_11509, n_11685);
  nand g26823 (n_11717, n_16232, n_16233);
  nand g26824 (n_15067, \data_stack_mem[8] [5], n_11716);
  nand g26825 (n_16234, n_12210, n_11748);
  or g26826 (n_16235, n_12210, n_11748);
  nand g26827 (n_11750, n_16234, n_16235);
  nand g26828 (n_11685, n_15042, n_15043);
  or g26829 (n_15046, \data_stack_mem[5] [7], n_11760);
  nand g26830 (n_11734, n_15012, n_15823);
  nand g26831 (n_16236, n_11699, n_11715);
  or g26832 (n_16237, n_11699, n_11715);
  nand g26833 (n_11716, n_16236, n_16237);
  nand g26834 (n_15007, n_15005, n_15006);
  nand g26835 (n_16238, n_11820, n_11823);
  or g26836 (n_16239, n_11820, n_11823);
  nand g26837 (n_11824, n_16238, n_16239);
  nand g26838 (n_11659, n_14946, n_14947);
  nand g26839 (n_11663, n_14964, n_14965);
  nand g26840 (n_11664, n_14970, n_14971);
  or g26842 (n_12210, n_15022, n_11515);
  nand g26843 (n_11661, n_14952, n_14953);
  nand g26844 (n_15823, n_11715, n_12207);
  nand g26845 (n_11657, n_14982, n_14983);
  or g26846 (n_15042, wc89, n_11506);
  not gc89 (wc89, n_12324);
  or g26847 (n_15005, \data_stack_mem[6] [6], n_11736);
  nand g26848 (n_15006, \data_stack_mem[6] [6], n_11736);
  nand g26849 (n_11662, n_14958, n_14959);
  nand g26850 (n_11660, n_14988, n_14989);
  nand g26851 (n_11658, n_14940, n_14941);
  nand g26852 (n_16240, n_11763, n_11771);
  or g26853 (n_16241, n_11763, n_11771);
  nand g26854 (n_11772, n_16240, n_16241);
  nand g26855 (n_16242, n_11780, n_11785);
  or g26856 (n_16243, n_11780, n_11785);
  nand g26857 (n_11786, n_16242, n_16243);
  nand g26858 (n_11760, n_15036, n_15037);
  nand g26859 (n_16244, n_11701, n_11714);
  or g26860 (n_16245, n_11701, n_11714);
  nand g26861 (n_11715, n_16244, n_16245);
  nand g26862 (n_15036, n_12312, n_11749);
  nand g26863 (n_11718, n_15030, n_15031);
  or g26864 (n_14983, n_11500, wc90);
  not gc90 (wc90, n_11656);
  nand g26865 (n_11736, n_14976, n_15820);
  or g26866 (n_14989, n_11544, wc91);
  not gc91 (wc91, n_11656);
  or g26867 (n_16246, wc92, n_11684);
  not gc92 (wc92, n_11683);
  or g26868 (n_16247, n_11683, wc93);
  not gc93 (wc93, n_11684);
  nand g26869 (n_12324, n_16246, n_16247);
  or g26870 (n_14970, n_11561, wc94);
  not gc94 (wc94, n_11656);
  nand g26871 (n_15013, n_12207, n_15012);
  or g26872 (n_11780, n_12258, wc95);
  not gc95 (wc95, n_15025);
  or g26873 (n_14965, n_11557, wc96);
  not gc96 (wc96, n_11656);
  or g26874 (n_14959, n_11553, wc97);
  not gc97 (wc97, n_11656);
  nand g26875 (n_15022, n_15020, n_15021);
  or g26876 (n_14953, n_11549, wc98);
  not gc98 (wc98, n_11656);
  or g26877 (n_14941, n_11536, wc99);
  not gc99 (wc99, n_11656);
  or g26878 (n_14947, n_11541, wc100);
  not gc100 (wc100, n_11656);
  nand g26879 (n_15030, n_12317, n_11682);
  nand g26883 (n_11683, n_16248, n_16249);
  nand g26884 (n_15037, \data_stack_mem[5] [6], n_11748);
  nand g26885 (n_15012, \data_stack_mem[7] [5], n_11698);
  nand g26887 (n_15021, \data_stack_mem[5] [6], n_11749);
  or g26888 (n_15020, \data_stack_mem[5] [6], n_11749);
  or g26890 (n_11701, n_14977, n_11513);
  nand g26892 (n_15820, n_12240, n_11714);
  nand g26893 (n_16250, n_11739, n_11747);
  or g26894 (n_16251, n_11739, n_11747);
  nand g26895 (n_11748, n_16250, n_16251);
  nand g26896 (n_16252, n_11666, n_11681);
  or g26897 (n_16253, n_11666, n_11681);
  nand g26898 (n_11682, n_16252, n_16253);
  nand g26899 (n_11698, n_14898, n_15814);
  nand g26900 (n_14977, n_12240, n_14976);
  nand g26901 (n_11749, n_14997, n_14998);
  nand g26902 (n_14935, n_14932, n_14933);
  or g26903 (n_14992, \data_stack_mem[4] [7], n_11762);
  nand g26906 (n_11823, n_11822, n_11821);
  nand g26907 (n_16256, n_12285, n_11712);
  or g26908 (n_16257, n_12285, n_11712);
  nand g26909 (n_11714, n_16256, n_16257);
  nand g26910 (n_16258, n_11781, n_11784);
  or g26911 (n_16259, n_11781, n_11784);
  nand g26912 (n_11785, n_16258, n_16259);
  nand g26913 (n_11762, n_14904, n_15817);
  nand g26914 (n_11630, n_14892, n_14893);
  or g26915 (n_12285, n_14818, n_11515);
  nand g26916 (n_11629, n_14886, n_14887);
  nand g26917 (n_11627, n_14874, n_14875);
  nand g26918 (n_16260, n_11765, n_11770);
  or g26919 (n_16261, n_11765, n_11770);
  nand g26920 (n_11771, n_16260, n_16261);
  nand g26921 (n_11625, n_14868, n_14869);
  or g26922 (n_11739, n_11516, n_14905);
  nand g26923 (n_14997, n_12286, n_11713);
  nand g26925 (n_11628, n_14880, n_14881);
  nand g26926 (n_11626, n_14916, n_14917);
  nand g26927 (n_14976, \data_stack_mem[6] [5], n_11700);
  nand g26928 (n_14933, n_11509, n_11652);
  nand g26929 (n_11623, n_14910, n_14911);
  nand g26930 (n_11624, n_14862, n_14863);
  nand g26931 (n_15814, n_12237, n_11681);
  or g26932 (n_14869, n_11541, wc101);
  not gc101 (wc101, n_11622);
  nand g26933 (n_14899, n_12237, n_14898);
  or g26934 (n_11781, n_12223, wc102);
  not gc102 (wc102, n_14920);
  nand g26935 (n_11652, n_14826, n_14827);
  nand g26936 (n_14998, \data_stack_mem[5] [5], n_11712);
  nand g26937 (n_14905, n_12271, n_14904);
  or g26938 (n_14887, n_11557, wc103);
  not gc103 (wc103, n_11622);
  or g26939 (n_14875, n_11549, wc104);
  not gc104 (wc104, n_11622);
  nand g26940 (n_16262, n_12252, n_11680);
  or g26941 (n_16263, n_12252, n_11680);
  nand g26942 (n_11681, n_16262, n_16263);
  or g26943 (n_14917, n_11544, wc105);
  not gc105 (wc105, n_11622);
  or g26944 (n_14863, n_11536, wc106);
  not gc106 (wc106, n_11622);
  or g26945 (n_14911, n_11500, wc107);
  not gc107 (wc107, n_11622);
  nand g26946 (n_15031, \data_stack_mem[8] [4], n_11684);
  nand g26947 (n_14818, n_14816, n_14817);
  or g26948 (n_14892, n_11561, wc108);
  not gc108 (wc108, n_11622);
  nand g26949 (n_15817, n_11747, n_12271);
  or g26950 (n_14881, n_11553, wc109);
  not gc109 (wc109, n_11622);
  nand g26951 (n_11700, n_14835, n_14836);
  or g26952 (n_12252, n_14713, n_11513);
  or g26953 (n_14826, n_14825, n_11506);
  nand g26955 (n_12223, n_11507, n_14830);
  nand g26956 (n_14898, \data_stack_mem[7] [4], n_11665);
  nand g26957 (n_14904, \data_stack_mem[4] [6], n_11738);
  nand g26958 (n_16264, n_11703, n_11711);
  or g26959 (n_16265, n_11703, n_11711);
  nand g26960 (n_11712, n_16264, n_16265);
  nand g26961 (n_14817, \data_stack_mem[5] [5], n_11713);
  or g26963 (n_14816, \data_stack_mem[5] [5], n_11713);
  nand g26964 (n_14835, n_12282, n_11667);
  nand g26965 (n_11684, n_14841, n_14842);
  nand g26966 (n_14713, n_14711, n_14712);
  nand g26967 (n_11713, n_14808, n_14809);
  nand g26968 (n_14836, \data_stack_mem[6] [4], n_11680);
  nand g26969 (n_11665, n_14703, n_15805);
  nand g26970 (n_11738, n_14772, n_15808);
  nand g26971 (n_14857, n_14854, n_14855);
  or g26972 (n_11703, n_11516, n_14773);
  nand g26973 (n_16266, n_11741, n_11746);
  or g26974 (n_16267, n_11741, n_11746);
  nand g26975 (n_11747, n_16266, n_16267);
  or g26977 (n_14830, \data_stack_mem[3] [7], n_11764);
  nand g26978 (n_14827, n_12338, n_11651);
  nand g26979 (n_14841, n_12321, n_11651);
  nand g26980 (n_15805, n_11650, n_12256);
  nand g26981 (n_14773, n_12229, n_14772);
  nand g26983 (n_15808, n_11711, n_12229);
  nand g26984 (n_16268, n_11634, n_11650);
  or g26985 (n_16269, n_11634, n_11650);
  nand g26986 (n_11651, n_16268, n_16269);
  or g26987 (n_14711, \data_stack_mem[6] [4], n_11667);
  nand g26988 (n_16270, n_11669, n_11679);
  or g26989 (n_16271, n_11669, n_11679);
  nand g26990 (n_11680, n_16270, n_16271);
  nand g26991 (n_11764, n_14778, n_15811);
  nand g26992 (n_14855, n_11509, n_11618);
  nand g26993 (n_14712, \data_stack_mem[6] [4], n_11667);
  nand g26994 (n_12338, n_11505, n_14800);
  nand g26995 (n_16272, n_11767, n_11769);
  or g26996 (n_16273, n_11767, n_11769);
  nand g26997 (n_11770, n_16272, n_16273);
  or g26998 (n_11821, n_11783, n_11782);
  nand g26999 (n_14808, n_12284, n_11668);
  or g27000 (n_16274, wc110, n_11783);
  not gc110 (wc110, n_11782);
  or g27001 (n_16275, n_11782, wc111);
  not gc111 (wc111, n_11783);
  nand g27002 (n_11784, n_16274, n_16275);
  nand g27003 (n_14809, \data_stack_mem[5] [4], n_11679);
  nand g27005 (n_14779, n_12272, n_14778);
  or g27006 (n_11669, n_14662, n_11515);
  nand g27007 (n_11618, n_14796, n_14797);
  nand g27008 (n_16276, n_11636, n_11649);
  or g27009 (n_16277, n_11636, n_11649);
  nand g27010 (n_11650, n_16276, n_16277);
  nand g27011 (n_11667, n_14673, n_15796);
  or g27012 (n_11782, n_12218, wc112);
  not gc112 (wc112, n_14803);
  nand g27013 (n_15811, n_11746, n_12272);
  or g27014 (n_14800, n_11506, n_11632);
  nand g27015 (n_14772, \data_stack_mem[4] [5], n_11702);
  nand g27016 (n_12218, n_11517, n_14716);
  nand g27017 (n_14842, \data_stack_mem[8] [3], n_11631);
  nand g27018 (n_11589, n_14784, n_14785);
  nand g27019 (n_11592, n_14790, n_14791);
  nand g27020 (n_11596, n_14766, n_14767);
  nand g27021 (n_11595, n_14760, n_14761);
  nand g27022 (n_15796, n_11649, n_12220);
  or g27023 (n_14796, wc113, n_11506);
  not gc113 (wc113, n_12334);
  or g27025 (n_11636, n_14674, n_11513);
  nand g27026 (n_11594, n_14754, n_14755);
  nand g27027 (n_14778, \data_stack_mem[3] [6], n_11740);
  nand g27028 (n_16278, n_11671, n_11678);
  or g27029 (n_16279, n_11671, n_11678);
  nand g27030 (n_11679, n_16278, n_16279);
  nand g27033 (n_11632, n_16280, n_16281);
  nand g27034 (n_11593, n_14748, n_14749);
  nand g27035 (n_14704, n_12256, n_14703);
  nand g27036 (n_14662, n_14660, n_14661);
  nand g27037 (n_16282, n_11705, n_11710);
  or g27038 (n_16283, n_11705, n_11710);
  nand g27039 (n_11711, n_16282, n_16283);
  nand g27040 (n_11702, n_14625, n_15778);
  nand g27041 (n_11591, n_14742, n_14743);
  nand g27042 (n_11590, n_14736, n_14737);
  nand g27043 (n_15778, n_12296, n_11678);
  or g27044 (n_14743, n_11541, wc114);
  not gc114 (wc114, n_11588);
  or g27045 (n_14785, n_11500, wc115);
  not gc115 (wc115, n_11588);
  nand g27046 (n_16284, n_11638, n_11648);
  or g27047 (n_16285, n_11638, n_11648);
  nand g27048 (n_11649, n_16284, n_16285);
  or g27049 (n_14761, n_11557, wc116);
  not gc116 (wc116, n_11588);
  or g27050 (n_11671, n_11516, n_14626);
  or g27051 (n_14755, n_11553, wc117);
  not gc117 (wc117, n_11588);
  nand g27052 (n_14674, n_12220, n_14673);
  nand g27053 (n_14703, \data_stack_mem[7] [3], n_11633);
  or g27054 (n_14749, n_11549, wc118);
  not gc118 (wc118, n_11588);
  or g27056 (n_16286, wc119, n_11617);
  not gc119 (wc119, n_11616);
  or g27057 (n_16287, n_11616, wc120);
  not gc120 (wc120, n_11617);
  nand g27058 (n_12334, n_16286, n_16287);
  or g27059 (n_14716, \data_stack_mem[2] [7], n_11766);
  nand g27060 (n_11740, n_14679, n_15799);
  or g27061 (n_14660, \data_stack_mem[5] [4], n_11668);
  nand g27062 (n_11631, n_14697, n_14698);
  nand g27063 (n_14661, \data_stack_mem[5] [4], n_11668);
  nand g27064 (n_16288, n_11743, n_11745);
  or g27065 (n_16289, n_11743, n_11745);
  nand g27066 (n_11746, n_16288, n_16289);
  or g27067 (n_14737, n_11536, wc121);
  not gc121 (wc121, n_11588);
  or g27068 (n_14791, n_11544, wc122);
  not gc122 (wc122, n_11588);
  or g27069 (n_14766, n_11561, wc123);
  not gc123 (wc123, n_11588);
  nand g27070 (n_14680, n_12179, n_14679);
  nand g27071 (n_11633, n_14640, n_15787);
  nand g27074 (n_14626, n_12296, n_14625);
  nand g27075 (n_11668, n_14646, n_15790);
  nand g27076 (n_14697, n_12322, n_11615);
  nand g27077 (n_11766, n_14685, n_15802);
  or g27078 (n_11638, n_14647, n_11515);
  or g27079 (n_11743, n_14686, wc124);
  not gc124 (wc124, n_11517);
  nand g27080 (n_11678, n_14667, n_14668);
  nand g27081 (n_15799, n_11710, n_12179);
  nand g27082 (n_14673, \data_stack_mem[6] [3], n_11635);
  nand g27085 (n_11616, n_16290, n_16291);
  nand g27086 (n_11635, n_14601, n_15775);
  nand g27087 (n_16292, n_11598, n_11614);
  or g27088 (n_16293, n_11598, n_11614);
  nand g27089 (n_11615, n_16292, n_16293);
  nand g27090 (n_14731, n_14728, n_14729);
  nand g27091 (n_14625, \data_stack_mem[4] [4], n_11670);
  nand g27092 (n_15790, n_11648, n_12221);
  or g27093 (n_14667, n_12287, n_11676);
  nand g27094 (n_15787, n_11614, n_12224);
  nand g27095 (n_14668, n_11676, n_12287);
  nand g27096 (n_14647, n_12221, n_14646);
  nand g27097 (n_14679, \data_stack_mem[3] [5], n_11704);
  nand g27098 (n_14686, n_12178, n_14685);
  nand g27099 (n_15802, n_12178, n_11745);
  nand g27100 (n_16294, n_11707, n_11709);
  or g27101 (n_16295, n_11707, n_11709);
  nand g27102 (n_11710, n_16294, n_16295);
  nand g27103 (n_14685, \data_stack_mem[2] [6], n_11742);
  nand g27104 (n_11670, n_14583, n_15769);
  nand g27105 (n_15775, n_12189, n_11613);
  nand g27106 (n_16296, n_11600, n_11613);
  or g27107 (n_16297, n_11600, n_11613);
  nand g27108 (n_11614, n_16296, n_16297);
  nand g27109 (n_16298, n_11640, n_11647);
  or g27110 (n_16299, n_11640, n_11647);
  nand g27111 (n_11648, n_16298, n_16299);
  nand g27112 (n_14646, \data_stack_mem[5] [3], n_11637);
  nand g27113 (n_14729, n_11509, n_11584);
  nand g27114 (n_11704, n_14652, n_15793);
  nand g27116 (n_11584, n_14691, n_14692);
  nand g27117 (n_11742, n_14631, n_15781);
  nand g27118 (n_11613, n_14616, n_14617);
  nand g27119 (n_16300, n_12236, \data_stack_mem[0] [7]);
  or g27120 (n_16301, n_12236, \data_stack_mem[0] [7]);
  nand g27121 (n_11769, n_16300, n_16301);
  nand g27122 (n_11637, n_14589, n_15772);
  or g27123 (n_11707, n_14632, wc125);
  not gc125 (wc125, n_11517);
  nand g27124 (n_15793, n_11676, n_12180);
  nand g27125 (n_14653, n_12180, n_14652);
  nand g27126 (n_15769, n_12283, n_11647);
  or g27127 (n_11640, n_11516, n_14584);
  nand g27128 (n_14584, n_12283, n_14583);
  or g27129 (n_14616, n_12314, n_11612);
  nand g27131 (n_14652, \data_stack_mem[3] [4], n_11677);
  nand g27132 (n_11647, n_14595, n_14596);
  or g27133 (n_14691, wc126, n_11506);
  not gc126 (wc126, n_12349);
  nand g27134 (n_14698, \data_stack_mem[8] [2], n_11617);
  nand g27135 (n_15772, n_12182, n_11612);
  or g27136 (n_12236, n_14443, wc127);
  not gc127 (wc127, n_11508);
  nand g27137 (n_11783, n_12353, n_11508);
  nand g27138 (n_14632, n_12214, n_14631);
  nand g27139 (n_15781, n_11709, n_12214);
  nand g27140 (n_14617, n_11612, n_12314);
  nand g27141 (n_11617, n_14635, n_15784);
  nand g27142 (n_14443, n_14441, n_14442);
  nand g27143 (n_11550, n_14538, n_14539);
  nand g27144 (n_12353, n_12126, n_14458);
  nand g27145 (n_11542, n_14532, n_14533);
  nand g27146 (n_14631, \data_stack_mem[2] [5], n_11706);
  nand g27147 (n_11537, n_14526, n_14527);
  nand g27148 (n_11677, n_14484, n_15763);
  nand g27149 (n_11554, n_14544, n_14545);
  or g27150 (n_14596, n_12299, wc128);
  not gc128 (wc128, n_11646);
  or g27151 (n_14595, wc129, n_11646);
  not gc129 (wc129, n_12299);
  nand g27152 (n_11558, n_14550, n_14551);
  nand g27153 (n_14583, \data_stack_mem[4] [3], n_11639);
  nand g27154 (n_11562, n_14556, n_14557);
  nand g27155 (n_11612, n_14514, n_14515);
  or g27156 (n_11600, n_14602, n_11513);
  nand g27157 (n_11531, n_14568, n_14569);
  nand g27158 (n_16302, n_11673, n_11675);
  or g27159 (n_16303, n_11673, n_11675);
  nand g27160 (n_11676, n_16302, n_16303);
  nand g27161 (n_16304, n_12242, \data_stack_mem[0] [6]);
  or g27162 (n_16305, n_12242, \data_stack_mem[0] [6]);
  nand g27163 (n_11745, n_16304, n_16305);
  or g27164 (n_16306, wc130, n_11583);
  not gc130 (wc130, n_11565);
  or g27165 (n_16307, n_11565, wc131);
  not gc131 (wc131, n_11583);
  nand g27166 (n_12349, n_16306, n_16307);
  nand g27167 (n_11545, n_14574, n_14575);
  nand g27168 (n_14641, n_12224, n_14640);
  nand g27170 (n_14640, \data_stack_mem[7] [2], n_11597);
  nand g27173 (n_12299, n_14493, n_14494);
  nand g27175 (n_15763, n_12293, n_11646);
  nand g27179 (n_14458, n_12352, n_11768);
  nand g27180 (n_14515, n_11610, n_12306);
  nand g27181 (n_11583, n_12257, n_14635);
  nand g27182 (n_11706, n_14562, n_15766);
  nand g27183 (n_14442, \data_stack_mem[1] [7], n_11768);
  or g27184 (n_14441, \data_stack_mem[1] [7], n_11768);
  or g27185 (n_14514, n_12306, n_11610);
  or g27186 (n_11673, n_14563, wc132);
  not gc132 (wc132, n_11517);
  or g27187 (n_15784, n_11565, wc133);
  not gc133 (wc133, n_12257);
  nand g27188 (n_11639, n_14454, n_15757);
  or g27190 (n_12314, n_14590, n_11515);
  nand g27191 (n_14602, n_12189, n_14601);
  or g27192 (n_12242, n_14413, wc134);
  not gc134 (wc134, n_11508);
  nand g27193 (n_14413, n_14411, n_14412);
  nand g27194 (n_15757, n_11610, n_12190);
  nand g27195 (n_16308, n_12204, \data_stack_mem[0] [5]);
  or g27196 (n_16309, n_12204, \data_stack_mem[0] [5]);
  nand g27197 (n_11709, n_16308, n_16309);
  nand g27198 (n_14635, \data_stack_mem[8] [1], n_11582);
  nand g27199 (n_14601, \data_stack_mem[6] [2], n_11599);
  nand g27201 (n_11646, n_14508, n_14509);
  nand g27202 (n_11597, n_14475, n_15760);
  nand g27203 (n_11768, n_12124, n_14434);
  nand g27204 (n_14590, n_12182, n_14589);
  nand g27205 (n_15766, n_12196, n_11675);
  or g27206 (n_12306, n_11516, n_14455);
  nand g27207 (n_11530, n_14520, n_14521);
  nand g27209 (n_14563, n_12196, n_14562);
  nand g27210 (n_11599, n_14402, n_15751);
  or g27211 (n_12058, n_13737, n_13738);
  or g27212 (n_12057, n_13689, n_13690);
  or g27213 (n_12066, n_14121, n_14122);
  nand g27214 (n_14562, \data_stack_mem[2] [4], n_11672);
  or g27215 (n_12063, n_13977, n_13978);
  nand g27216 (n_14589, \data_stack_mem[5] [2], n_11601);
  or g27217 (n_12059, n_13785, n_13786);
  nand g27218 (n_14434, n_12328, n_11744);
  or g27219 (n_12056, n_13641, n_13642);
  nand g27220 (n_16310, n_11603, n_11609);
  or g27221 (n_16311, n_11603, n_11609);
  nand g27222 (n_11610, n_16310, n_16311);
  or g27223 (n_12065, n_14073, n_14074);
  or g27224 (n_12053, n_13497, n_13498);
  or g27225 (n_12060, n_13833, n_13834);
  nand g27226 (n_14484, \data_stack_mem[3] [3], n_11641);
  or g27227 (n_12069, n_14265, n_14266);
  or g27228 (n_12055, n_13593, n_13594);
  or g27229 (n_12067, n_14169, n_14170);
  nand g27230 (n_16312, n_11567, n_11581);
  or g27231 (n_16313, n_11567, n_11581);
  nand g27232 (n_11582, n_16312, n_16313);
  or g27233 (n_12062, n_13929, n_13930);
  nand g27234 (n_14509, n_11645, n_12289);
  nand g27235 (n_14455, n_12190, n_14454);
  or g27236 (n_14508, n_12289, n_11645);
  or g27237 (n_12064, n_14025, n_14026);
  nand g27238 (n_14520, n_12366, n_11509);
  or g27240 (n_14492, wc135, n_11641);
  not gc135 (wc135, \data_stack_mem[3] [3]);
  or g27241 (n_12204, n_14386, wc136);
  not gc136 (wc136, n_11508);
  or g27242 (n_12061, n_13881, n_13882);
  nand g27243 (n_14412, \data_stack_mem[1] [6], n_11744);
  or g27244 (n_12054, n_13545, n_13546);
  or g27245 (n_14411, \data_stack_mem[1] [6], n_11744);
  nand g27246 (n_15760, n_11581, n_12259);
  or g27247 (n_12068, n_14217, n_14218);
  or g27249 (n_13738, n_13735, n_13736);
  or g27250 (n_13690, n_13687, n_13688);
  nand g27252 (n_14386, n_14384, n_14385);
  or g27253 (n_13786, n_13783, n_13784);
  or g27254 (n_13642, n_13639, n_13640);
  nand g27255 (n_16314, n_12219, n_11580);
  or g27256 (n_16315, n_12219, n_11580);
  nand g27257 (n_11581, n_16314, n_16315);
  or g27258 (n_14074, n_14071, n_14072);
  or g27259 (n_13834, n_13831, n_13832);
  nand g27260 (n_14454, \data_stack_mem[4] [2], n_11611);
  or g27261 (n_13594, n_13591, n_13592);
  or g27262 (n_13882, n_13879, n_13880);
  or g27263 (n_13978, n_13975, n_13976);
  or g27264 (n_12009, n_14307, n_14308);
  or g27265 (n_12289, n_14449, wc137);
  not gc137 (wc137, n_11517);
  or g27266 (n_14170, n_14167, n_14168);
  nand g27267 (n_15751, n_12316, n_11580);
  or g27268 (n_13546, n_13543, n_13544);
  nand g27269 (n_11672, n_14448, n_15754);
  nand g27270 (n_11601, n_14394, n_15748);
  nand g27271 (n_11641, n_14316, n_15739);
  or g27272 (n_14266, n_14263, n_14264);
  or g27273 (n_14026, n_14023, n_14024);
  or g27274 (n_15345, n_15342, wc138);
  not gc138 (wc138, n_12153);
  or g27275 (n_14122, n_14119, n_14120);
  nand g27276 (n_16316, n_12254, \data_stack_mem[0] [4]);
  or g27277 (n_16317, n_12254, \data_stack_mem[0] [4]);
  nand g27278 (n_11675, n_16316, n_16317);
  or g27279 (n_13498, n_13495, n_13496);
  nand g27280 (n_11744, n_12122, n_14389);
  or g27281 (n_14218, n_14215, n_14216);
  or g27282 (n_13930, n_13927, n_13928);
  or g27290 (n_15081, n_11688, n_15078);
  nand g27291 (n_14449, n_12216, n_14448);
  or g27292 (n_14856, n_11621, n_14853);
  nand g27293 (n_15754, n_11645, n_12216);
  nand g27295 (n_15739, n_12297, n_11609);
  or g27296 (n_15342, n_15340, n_15341);
  or g27297 (n_12254, n_13036, wc139);
  not gc139 (wc139, n_11508);
  nand g27300 (n_14470, n_11522, n_14468);
  or g27301 (n_15261, n_11756, n_15258);
  nand g27302 (n_16318, n_11570, n_11579);
  or g27303 (n_16319, n_11570, n_11579);
  nand g27304 (n_11580, n_16318, n_16319);
  or g27306 (n_14308, n_14305, n_14306);
  or g27307 (n_14730, n_11587, n_14727);
  or g27308 (n_14307, n_14303, n_14304);
  or g27311 (n_15177, n_11722, n_15174);
  or g27314 (n_14934, n_11655, n_14931);
  or g27315 (n_14384, \data_stack_mem[1] [5], n_11708);
  nand g27318 (n_14385, \data_stack_mem[1] [5], n_11708);
  nand g27319 (n_14317, n_12297, n_14316);
  nand g27320 (n_11611, n_14328, n_15745);
  nand g27321 (n_15748, n_11579, n_12225);
  nand g27323 (n_14389, n_12327, n_11708);
  nand g27324 (n_11994, n_13317, n_13318);
  nand g27325 (n_13540, n_13531, n_13532);
  nand g27326 (n_11972, n_14334, n_14335);
  nand g27327 (n_11993, n_13311, n_13312);
  nand g27328 (n_14020, n_14011, n_14012);
  nand g27329 (n_13543, n_13537, n_13538);
  nand g27330 (n_11990, n_13305, n_13306);
  nand g27331 (n_15258, n_12311, n_12310);
  or g27332 (n_13545, n_13541, n_13542);
  nand g27333 (n_11989, n_13299, n_13300);
  nand g27334 (n_16320, n_11572, n_11578);
  or g27335 (n_16321, n_11572, n_11578);
  nand g27336 (n_11579, n_16320, n_16321);
  nand g27337 (n_11977, n_14364, n_14365);
  nand g27338 (n_11988, n_13293, n_13294);
  nand g27339 (n_11995, n_13323, n_13324);
  nand g27340 (n_14023, n_14017, n_14018);
  nand g27341 (n_11987, n_13287, n_13288);
  nand g27342 (n_14853, n_12336, n_12335);
  nand g27343 (n_11996, n_13329, n_13330);
  nand g27344 (n_11986, n_13281, n_13282);
  or g27345 (n_14025, n_14021, n_14022);
  nand g27346 (n_13876, n_13867, n_13868);
  nand g27347 (n_11985, n_13275, n_13276);
  nand g27348 (n_11997, n_13335, n_13336);
  nand g27349 (n_14164, n_14155, n_14156);
  nand g27350 (n_11984, n_13269, n_13270);
  nand g27351 (n_13684, n_13675, n_13676);
  nand g27352 (n_11998, n_13341, n_13342);
  nand g27353 (n_11983, n_13263, n_13264);
  nand g27354 (n_11897, n_13407, n_13408);
  nand g27355 (n_12035, n_12984, n_12985);
  nand g27356 (n_11921, n_13257, n_13258);
  nand g27357 (n_14931, n_12340, n_12339);
  nand g27358 (n_11999, n_13347, n_13348);
  nand g27359 (n_11920, n_13251, n_13252);
  nand g27360 (n_11973, n_14340, n_14341);
  nand g27361 (n_13879, n_13873, n_13874);
  nand g27362 (n_11919, n_13245, n_13246);
  nand g27363 (n_12000, n_13353, n_13354);
  nand g27364 (n_13687, n_13681, n_13682);
  nand g27365 (n_11918, n_13239, n_13240);
  or g27366 (n_13689, n_13685, n_13686);
  or g27367 (n_13881, n_13877, n_13878);
  nand g27368 (n_11917, n_13233, n_13234);
  nand g27369 (n_12052, n_12966, n_12967);
  nand g27370 (n_14260, n_14251, n_14252);
  nand g27371 (n_11916, n_13227, n_13228);
  nand g27372 (n_14167, n_14161, n_14162);
  nand g27373 (n_12051, n_12960, n_12961);
  nand g27374 (n_11915, n_13221, n_13222);
  nand g27375 (n_11708, n_12120, n_13096);
  or g27376 (n_12219, n_14404, n_11513);
  nand g27377 (n_11914, n_13215, n_13216);
  nand g27378 (n_12050, n_12954, n_12955);
  nand g27379 (n_12039, n_12900, n_12901);
  nand g27380 (n_14263, n_14257, n_14258);
  nand g27381 (n_12049, n_12948, n_12949);
  or g27382 (n_14169, n_14165, n_14166);
  nand g27383 (n_13492, n_13483, n_13484);
  nand g27384 (n_12048, n_12942, n_12943);
  or g27385 (n_14468, n_14467, n_11506);
  nand g27386 (n_14068, n_14059, n_14060);
  nand g27387 (n_12047, n_12936, n_12937);
  nand g27388 (n_13732, n_13723, n_13724);
  nand g27389 (n_11898, n_13413, n_13414);
  nand g27390 (n_12046, n_12930, n_12931);
  or g27391 (n_14265, n_14261, n_14262);
  nand g27392 (n_13924, n_13915, n_13916);
  nand g27393 (n_12045, n_12924, n_12925);
  nand g27394 (n_11899, n_13419, n_13420);
  nand g27395 (n_13735, n_13729, n_13730);
  or g27396 (n_13737, n_13733, n_13734);
  nand g27397 (n_12042, n_12918, n_12919);
  nand g27398 (n_11974, n_14346, n_14347);
  nand g27399 (n_11900, n_13425, n_13426);
  nand g27400 (n_12041, n_12912, n_12913);
  nand g27401 (n_15174, n_12320, n_12319);
  nand g27402 (n_14071, n_14065, n_14066);
  nand g27403 (n_12040, n_12906, n_12907);
  nand g27404 (n_11880, n_13161, n_13162);
  nand g27405 (n_13927, n_13921, n_13922);
  nand g27406 (n_13588, n_13579, n_13580);
  nand g27407 (n_11879, n_13155, n_13156);
  nand g27408 (n_15078, n_12326, n_12325);
  or g27409 (n_13929, n_13925, n_13926);
  nand g27410 (n_11878, n_13149, n_13150);
  or g27411 (n_14073, n_14069, n_14070);
  nand g27412 (n_12037, n_12894, n_12895);
  nand g27413 (n_11877, n_13143, n_13144);
  nand g27414 (n_13036, n_13034, n_13035);
  nand g27415 (n_11978, n_14370, n_14371);
  nand g27416 (n_11876, n_13137, n_13138);
  nand g27417 (n_12036, n_12888, n_12889);
  nand g27418 (n_16322, n_11605, n_11608);
  or g27419 (n_16323, n_11605, n_11608);
  nand g27420 (n_11609, n_16322, n_16323);
  nand g27421 (n_11875, n_13131, n_13132);
  nand g27422 (n_15745, n_11578, n_12238);
  nand g27423 (n_11979, n_14376, n_14377);
  nand g27424 (n_11874, n_13125, n_13126);
  nand g27425 (n_13780, n_13771, n_13772);
  nand g27426 (n_14316, \data_stack_mem[3] [2], n_11602);
  nand g27427 (n_11873, n_13119, n_13120);
  nand g27428 (n_13783, n_13777, n_13778);
  or g27429 (n_13785, n_13781, n_13782);
  nand g27430 (n_14212, n_14203, n_14204);
  nand g27431 (n_11901, n_13431, n_13432);
  nand g27432 (n_13495, n_13489, n_13490);
  or g27433 (n_13497, n_13493, n_13494);
  nand g27434 (n_11902, n_13437, n_13438);
  nand g27435 (n_14303, n_14295, n_14296);
  nand g27436 (n_14116, n_14107, n_14108);
  nand g27437 (n_11903, n_13443, n_13444);
  nand g27438 (n_13972, n_13963, n_13964);
  nand g27439 (n_11975, n_14352, n_14353);
  nand g27440 (n_14727, n_12351, n_12350);
  nand g27441 (n_13591, n_13585, n_13586);
  or g27442 (n_13593, n_13589, n_13590);
  nand g27443 (n_14215, n_14209, n_14210);
  nand g27444 (n_13975, n_13969, n_13970);
  or g27445 (n_15341, wc140, n_11813);
  not gc140 (wc140, n_12200);
  or g27446 (n_13977, n_13973, n_13974);
  nand g27447 (n_14119, n_14113, n_14114);
  or g27448 (n_14121, n_14117, n_14118);
  or g27449 (n_14217, n_14213, n_14214);
  nand g27450 (n_13828, n_13819, n_13820);
  nand g27451 (n_14305, n_14299, n_14300);
  nand g27452 (n_14448, \data_stack_mem[2] [3], n_11642);
  nand g27453 (n_13636, n_13627, n_13628);
  nand g27454 (n_13831, n_13825, n_13826);
  or g27455 (n_13833, n_13829, n_13830);
  nand g27456 (n_11904, n_13449, n_13450);
  nand g27457 (n_13639, n_13633, n_13634);
  or g27458 (n_13641, n_13637, n_13638);
  nand g27459 (n_11976, n_14358, n_14359);
  nand g27460 (n_12038, n_13026, n_13027);
  nand g27461 (n_14476, n_12259, n_14475);
  nand g27462 (n_13426, \data_stack_mem[0] [3], n_11895);
  nand g27463 (n_16324, n_11644, \data_stack_mem[0] [3]);
  or g27464 (n_16325, n_11644, \data_stack_mem[0] [3]);
  nand g27465 (n_11645, n_16324, n_16325);
  nand g27466 (n_13318, \data_stack_mem[7] [1], n_11991);
  nand g27467 (n_14377, \data_stack_mem[5] [3], n_11971);
  nand g27468 (n_13312, \data_stack_mem[7] [7], n_11991);
  nand g27469 (n_14371, \data_stack_mem[5] [0], n_11971);
  nand g27470 (n_13306, \data_stack_mem[6] [7], n_11982);
  or g27471 (n_13633, wc141, n_12006);
  not gc141 (wc141, \out_fifo[0][1] [1]);
  nand g27472 (n_13300, \data_stack_mem[6] [3], n_11982);
  or g27473 (n_14011, wc142, n_12073);
  not gc142 (wc142, \out_fifo[4][0] [2]);
  nand g27474 (n_13294, \data_stack_mem[6] [2], n_11982);
  nand g27475 (n_13974, n_13967, n_13968);
  nand g27476 (n_13288, \data_stack_mem[6] [1], n_11982);
  nand g27477 (n_13973, n_13965, n_13966);
  nand g27478 (n_13282, \data_stack_mem[6] [6], n_11982);
  nand g27479 (n_13354, \data_stack_mem[7] [2], n_11991);
  nand g27480 (n_13276, \data_stack_mem[6] [5], n_11982);
  nand g27481 (n_13444, \data_stack_mem[0] [6], n_11895);
  nand g27482 (n_13270, \data_stack_mem[6] [4], n_11982);
  or g27483 (n_13969, wc143, n_12006);
  not gc143 (wc143, \out_fifo[0][0] [3]);
  nand g27484 (n_13264, \data_stack_mem[6] [0], n_11982);
  nand g27485 (n_12340, n_11564, n_12754);
  nand g27486 (n_13258, \data_stack_mem[2] [7], n_11913);
  nand g27487 (n_11487, n_13359, n_13360);
  nand g27488 (n_13252, \data_stack_mem[2] [0], n_11913);
  nand g27489 (n_13438, \data_stack_mem[0] [5], n_11895);
  nand g27490 (n_13246, \data_stack_mem[2] [6], n_11913);
  or g27491 (n_11570, n_14395, n_11515);
  nand g27492 (n_13240, \data_stack_mem[2] [4], n_11913);
  or g27493 (n_13963, wc144, n_12073);
  not gc144 (wc144, \out_fifo[4][0] [3]);
  nand g27494 (n_13234, \data_stack_mem[2] [5], n_11913);
  nand g27495 (n_13926, n_13919, n_13920);
  nand g27496 (n_13228, \data_stack_mem[2] [3], n_11913);
  nand g27497 (n_11492, n_13389, n_13390);
  nand g27498 (n_13222, \data_stack_mem[2] [2], n_11913);
  or g27499 (n_13627, wc145, n_12073);
  not gc145 (wc145, \out_fifo[4][1] [1]);
  nand g27500 (n_13216, \data_stack_mem[2] [1], n_11913);
  nand g27501 (n_13590, n_13583, n_13584);
  nand g27502 (n_11892, n_13209, n_13210);
  nand g27503 (n_14365, \data_stack_mem[5] [2], n_11971);
  or g27504 (n_13921, wc146, n_12006);
  not gc146 (wc146, \out_fifo[0][0] [4]);
  nand g27505 (n_11891, n_13203, n_13204);
  nand g27506 (n_14359, \data_stack_mem[5] [5], n_11971);
  nand g27507 (n_13589, n_13581, n_13582);
  nand g27508 (n_11890, n_13197, n_13198);
  nand g27509 (n_14353, \data_stack_mem[5] [6], n_11971);
  nand g27510 (n_11642, n_14322, n_15742);
  nand g27511 (n_11889, n_13191, n_13192);
  or g27512 (n_13483, wc147, n_12073);
  not gc147 (wc147, \out_fifo[4][1] [3]);
  nand g27513 (n_11488, n_13365, n_13366);
  nand g27514 (n_11888, n_13185, n_13186);
  or g27515 (n_13034, \data_stack_mem[1] [4], n_11674);
  or g27516 (n_13915, wc148, n_12073);
  not gc148 (wc148, \out_fifo[4][0] [4]);
  nand g27517 (n_11887, n_13179, n_13180);
  nand g27518 (n_13035, \data_stack_mem[1] [4], n_11674);
  nand g27519 (n_13878, n_13871, n_13872);
  nand g27520 (n_11886, n_13173, n_13174);
  nand g27521 (n_14347, \data_stack_mem[5] [4], n_11971);
  nand g27522 (n_13877, n_13869, n_13870);
  nand g27523 (n_11885, n_13167, n_13168);
  nand g27524 (n_14341, \data_stack_mem[5] [7], n_11971);
  nand g27525 (n_12326, n_11564, n_12748);
  nand g27526 (n_13162, \data_stack_mem[3] [6], n_11872);
  nand g27527 (n_14335, \data_stack_mem[5] [1], n_11971);
  nand g27528 (n_13156, \data_stack_mem[3] [3], n_11872);
  nand g27529 (n_14306, n_14301, n_14302);
  nand g27530 (n_13150, \data_stack_mem[3] [2], n_11872);
  nand g27531 (n_14304, n_14297, n_14298);
  nand g27532 (n_13144, \data_stack_mem[3] [1], n_11872);
  nand g27533 (n_11494, n_13401, n_13402);
  nand g27534 (n_13138, \data_stack_mem[3] [5], n_11872);
  or g27535 (n_13873, wc149, n_12006);
  not gc149 (wc149, \out_fifo[0][0] [7]);
  nand g27536 (n_13132, \data_stack_mem[3] [0], n_11872);
  or g27537 (n_14300, wc150, n_12006);
  not gc150 (wc150, \out_fifo[0][0] [0]);
  nand g27538 (n_13126, \data_stack_mem[3] [4], n_11872);
  nand g27539 (n_13432, \data_stack_mem[0] [4], n_11895);
  nand g27540 (n_13120, \data_stack_mem[3] [7], n_11872);
  nand g27541 (n_11489, n_13371, n_13372);
  or g27542 (n_13585, wc151, n_12006);
  not gc151 (wc151, \out_fifo[0][2] [9]);
  nand g27543 (n_13420, \data_stack_mem[0] [2], n_11895);
  or g27544 (n_13867, wc152, n_12073);
  not gc152 (wc152, \out_fifo[4][0] [7]);
  or g27545 (n_14295, wc153, n_12073);
  not gc153 (wc153, \out_fifo[4][0] [0]);
  nand g27546 (n_14262, n_14255, n_14256);
  nand g27547 (n_14261, n_14253, n_14254);
  nand g27548 (n_13830, n_13823, n_13824);
  nand g27549 (n_13829, n_13821, n_13822);
  nand g27550 (n_11578, n_13092, n_13093);
  nand g27551 (n_11490, n_13377, n_13378);
  or g27552 (n_14257, wc154, n_12006);
  not gc154 (wc154, \out_fifo[0][2] [1]);
  or g27553 (n_13825, wc155, n_12006);
  not gc155 (wc155, \out_fifo[0][0] [5]);
  nand g27554 (n_13450, \data_stack_mem[0] [7], n_11895);
  or g27555 (n_11605, n_14323, wc156);
  not gc156 (wc156, n_11517);
  nand g27556 (n_12336, n_11564, n_12751);
  nand g27557 (n_11491, n_13383, n_13384);
  or g27558 (n_13819, wc157, n_12073);
  not gc157 (wc157, \out_fifo[4][0] [5]);
  or g27559 (n_14251, wc158, n_12073);
  not gc158 (wc158, \out_fifo[4][2] [1]);
  nand g27560 (n_13782, n_13775, n_13776);
  nand g27561 (n_14214, n_14207, n_14208);
  nand g27562 (n_14213, n_14205, n_14206);
  nand g27563 (n_13781, n_13773, n_13774);
  nand g27564 (n_13408, \data_stack_mem[0] [0], n_11895);
  or g27565 (n_13579, wc159, n_12073);
  not gc159 (wc159, \out_fifo[4][2] [9]);
  or g27566 (n_13777, wc160, n_12006);
  not gc160 (wc160, \out_fifo[0][0] [6]);
  or g27567 (n_14209, wc161, n_12006);
  not gc161 (wc161, \out_fifo[0][1] [4]);
  nand g27568 (n_13542, n_13535, n_13536);
  nand g27569 (n_13541, n_13533, n_13534);
  nand g27570 (n_13414, \data_stack_mem[0] [1], n_11895);
  nand g27571 (n_11493, n_13395, n_13396);
  nand g27572 (n_12320, n_11564, n_12745);
  or g27573 (n_14203, wc162, n_12073);
  not gc162 (wc162, \out_fifo[4][1] [4]);
  or g27574 (n_13027, n_12034, n_11544);
  nand g27575 (n_13096, n_12323, n_11674);
  nand g27576 (n_11964, n_13020, n_13021);
  nand g27577 (n_14166, n_14159, n_14160);
  or g27578 (n_13771, wc163, n_12073);
  not gc163 (wc163, \out_fifo[4][0] [6]);
  nand g27579 (n_11963, n_13014, n_13015);
  nand g27580 (n_13734, n_13727, n_13728);
  nand g27581 (n_14165, n_14157, n_14158);
  nand g27582 (n_11962, n_13008, n_13009);
  nand g27583 (n_13733, n_13725, n_13726);
  nand g27584 (n_12200, n_12730, n_11564);
  nand g27585 (n_11961, n_13002, n_13003);
  or g27586 (n_13537, wc164, n_12006);
  not gc164 (wc164, \out_fifo[0][1] [2]);
  or g27587 (n_13729, wc165, n_12006);
  not gc165 (wc165, \out_fifo[0][2] [8]);
  nand g27588 (n_11960, n_12996, n_12997);
  or g27589 (n_13489, wc166, n_12006);
  not gc166 (wc166, \out_fifo[0][1] [3]);
  or g27590 (n_14161, wc167, n_12006);
  not gc167 (wc167, \out_fifo[0][2] [0]);
  nand g27591 (n_11959, n_12990, n_12991);
  nand g27592 (n_12351, n_11564, n_12757);
  nand g27593 (n_11602, n_12831, n_15736);
  or g27594 (n_12985, n_12034, n_11500);
  nand g27595 (n_12311, n_11564, n_12742);
  nand g27596 (n_11956, n_12978, n_12979);
  nand g27597 (n_13925, n_13917, n_13918);
  nand g27598 (n_11955, n_12972, n_12973);
  or g27599 (n_13531, wc168, n_12073);
  not gc168 (wc168, \out_fifo[4][1] [2]);
  nand g27600 (n_12967, \data_stack_mem[4] [0], n_12043);
  or g27601 (n_14155, wc169, n_12073);
  not gc169 (wc169, \out_fifo[4][2] [0]);
  nand g27602 (n_12961, \data_stack_mem[4] [1], n_12043);
  nand g27603 (n_14118, n_14111, n_14112);
  nand g27604 (n_12955, \data_stack_mem[4] [2], n_12043);
  nand g27605 (n_14117, n_14109, n_14110);
  nand g27606 (n_12949, \data_stack_mem[4] [4], n_12043);
  or g27607 (n_13723, wc170, n_12073);
  not gc170 (wc170, \out_fifo[4][2] [8]);
  nand g27608 (n_12943, \data_stack_mem[4] [3], n_12043);
  nand g27609 (n_13686, n_13679, n_13680);
  nand g27610 (n_12937, \data_stack_mem[4] [6], n_12043);
  or g27611 (n_14113, wc171, n_12006);
  not gc171 (wc171, \out_fifo[0][1] [0]);
  nand g27612 (n_12931, \data_stack_mem[4] [5], n_12043);
  nand g27613 (n_13685, n_13677, n_13678);
  nand g27614 (n_12925, \data_stack_mem[4] [7], n_12043);
  nand g27615 (n_13324, \data_stack_mem[7] [5], n_11991);
  nand g27616 (n_13494, n_13487, n_13488);
  or g27617 (n_14475, wc172, n_11566);
  not gc172 (wc172, \data_stack_mem[7] [1]);
  or g27618 (n_12918, n_11561, n_12034);
  or g27619 (n_12913, n_11557, n_12034);
  or g27620 (n_13681, wc173, n_12006);
  not gc173 (wc173, \out_fifo[0][0] [8]);
  or g27621 (n_12907, n_11553, n_12034);
  or g27622 (n_14107, wc174, n_12073);
  not gc174 (wc174, \out_fifo[4][1] [0]);
  nand g27623 (n_14070, n_14063, n_14064);
  or g27624 (n_12901, n_11549, n_12034);
  nand g27625 (n_14069, n_14061, n_14062);
  or g27626 (n_12895, n_11541, n_12034);
  nand g27627 (n_13330, \data_stack_mem[7] [6], n_11991);
  or g27628 (n_12889, n_11536, n_12034);
  nand g27629 (n_13493, n_13485, n_13486);
  nand g27630 (n_13336, \data_stack_mem[7] [0], n_11991);
  or g27631 (n_14065, wc175, n_12006);
  not gc175 (wc175, \out_fifo[0][0] [1]);
  nand g27632 (n_14469, n_12365, n_11529);
  nand g27633 (n_13342, \data_stack_mem[7] [4], n_11991);
  or g27634 (n_13675, wc176, n_12073);
  not gc176 (wc176, \out_fifo[4][0] [8]);
  or g27635 (n_14467, wc177, n_11529);
  not gc177 (wc177, \data_stack_mem[8] [0]);
  or g27636 (n_14059, wc178, n_12073);
  not gc178 (wc178, \out_fifo[4][0] [1]);
  nand g27637 (n_14022, n_14015, n_14016);
  nand g27638 (n_14021, n_14013, n_14014);
  nand g27639 (n_13638, n_13631, n_13632);
  nand g27640 (n_13637, n_13629, n_13630);
  or g27641 (n_14017, wc179, n_12006);
  not gc179 (wc179, \out_fifo[0][0] [2]);
  nand g27642 (n_13348, \data_stack_mem[7] [3], n_11991);
  nand g27643 (n_14404, n_12316, n_14402);
  or g27644 (n_11644, n_12823, wc180);
  not gc180 (wc180, n_11508);
  or g27645 (n_13305, wc181, n_11980);
  not gc181 (wc181, sh_reg_in[7]);
  or g27646 (n_13299, wc182, n_11980);
  not gc182 (wc182, sh_reg_in[3]);
  or g27647 (n_13293, wc183, n_11980);
  not gc183 (wc183, sh_reg_in[2]);
  or g27648 (n_13287, wc184, n_11980);
  not gc184 (wc184, sh_reg_in[1]);
  or g27649 (n_13281, wc185, n_11980);
  not gc185 (wc185, sh_reg_in[6]);
  or g27650 (n_13275, wc186, n_11980);
  not gc186 (wc186, sh_reg_in[5]);
  or g27651 (n_13269, wc187, n_11980);
  not gc187 (wc187, sh_reg_in[4]);
  or g27652 (n_13263, wc188, n_11980);
  not gc188 (wc188, sh_reg_in[0]);
  or g27653 (n_13257, wc189, n_11912);
  not gc189 (wc189, sh_reg_in[7]);
  or g27654 (n_13251, wc190, n_11912);
  not gc190 (wc190, sh_reg_in[0]);
  or g27655 (n_13245, wc191, n_11912);
  not gc191 (wc191, sh_reg_in[6]);
  or g27656 (n_13239, wc192, n_11912);
  not gc192 (wc192, sh_reg_in[4]);
  or g27657 (n_13233, wc193, n_11912);
  not gc193 (wc193, sh_reg_in[5]);
  or g27658 (n_13227, wc194, n_11912);
  not gc194 (wc194, sh_reg_in[3]);
  or g27659 (n_13221, wc195, n_11912);
  not gc195 (wc195, sh_reg_in[2]);
  or g27660 (n_13215, wc196, n_11912);
  not gc196 (wc196, sh_reg_in[1]);
  nand g27661 (n_13209, \data_stack_mem[1] [0], n_11884);
  nand g27662 (n_13203, \data_stack_mem[1] [1], n_11884);
  nand g27663 (n_13197, \data_stack_mem[1] [2], n_11884);
  nand g27664 (n_11674, n_12822, n_15733);
  nand g27665 (n_13191, \data_stack_mem[1] [3], n_11884);
  nand g27666 (n_13185, \data_stack_mem[1] [4], n_11884);
  nand g27667 (n_13179, \data_stack_mem[1] [5], n_11884);
  nand g27668 (n_13173, \data_stack_mem[1] [6], n_11884);
  nand g27669 (n_13167, \data_stack_mem[1] [7], n_11884);
  or g27670 (n_14302, wc197, n_12008);
  not gc197 (wc197, \out_fifo[2][0] [0]);
  or g27671 (n_14301, wc198, n_12007);
  not gc198 (wc198, \out_fifo[1][0] [0]);
  or g27672 (n_14299, wc199, n_12005);
  not gc199 (wc199, \out_fifo[3][0] [0]);
  or g27673 (n_14298, wc200, n_12070);
  not gc200 (wc200, \out_fifo[5][0] [0]);
  nand g27674 (n_11971, n_11485, n_13108);
  or g27675 (n_14297, wc201, n_12071);
  not gc201 (wc201, \out_fifo[6][0] [0]);
  or g27676 (n_14296, wc202, n_12072);
  not gc202 (wc202, \out_fifo[7][0] [0]);
  nand g27677 (n_11911, n_13086, n_13087);
  or g27678 (n_14259, wc203, n_12008);
  not gc203 (wc203, \out_fifo[2][2] [1]);
  or g27679 (n_14258, wc204, n_12007);
  not gc204 (wc204, \out_fifo[1][2] [1]);
  nand g27680 (n_11910, n_13080, n_13081);
  or g27681 (n_14256, wc205, n_12005);
  not gc205 (wc205, \out_fifo[3][2] [1]);
  nand g27682 (n_11958, n_13074, n_13075);
  or g27683 (n_14254, wc206, n_12070);
  not gc206 (wc206, \out_fifo[5][2] [1]);
  or g27684 (n_14253, wc207, n_12071);
  not gc207 (wc207, \out_fifo[6][2] [1]);
  nand g27685 (n_12030, n_13068, n_13069);
  or g27686 (n_14252, wc208, n_12072);
  not gc208 (wc208, \out_fifo[7][2] [1]);
  nand g27687 (n_12033, n_13062, n_13063);
  nand g27688 (n_12031, n_13056, n_13057);
  or g27689 (n_14211, wc209, n_12008);
  not gc209 (wc209, \out_fifo[2][1] [4]);
  or g27690 (n_14210, wc210, n_12007);
  not gc210 (wc210, \out_fifo[1][1] [4]);
  nand g27691 (n_11909, n_13050, n_13051);
  or g27692 (n_14208, wc211, n_12005);
  not gc211 (wc211, \out_fifo[3][1] [4]);
  nand g27693 (n_12032, n_13044, n_13045);
  or g27694 (n_14206, wc212, n_12070);
  not gc212 (wc212, \out_fifo[5][1] [4]);
  or g27695 (n_14205, wc213, n_12071);
  not gc213 (wc213, \out_fifo[6][1] [4]);
  or g27696 (n_14204, wc214, n_12072);
  not gc214 (wc214, \out_fifo[7][1] [4]);
  or g27697 (n_13020, n_11511, n_11561);
  or g27698 (n_13015, n_11511, n_11557);
  or g27699 (n_13009, n_11511, n_11553);
  or g27700 (n_14163, wc215, n_12008);
  not gc215 (wc215, \out_fifo[2][2] [0]);
  or g27701 (n_13003, n_11511, n_11549);
  or g27702 (n_14162, wc216, n_12007);
  not gc216 (wc216, \out_fifo[1][2] [0]);
  or g27703 (n_12997, n_11511, n_11541);
  or g27704 (n_12991, n_11511, n_11536);
  or g27705 (n_14160, wc217, n_12005);
  not gc217 (wc217, \out_fifo[3][2] [0]);
  or g27706 (n_14158, wc218, n_12070);
  not gc218 (wc218, \out_fifo[5][2] [0]);
  or g27707 (n_12979, n_11511, n_11544);
  or g27708 (n_14157, wc219, n_12071);
  not gc219 (wc219, \out_fifo[6][2] [0]);
  or g27709 (n_12973, n_11511, n_11500);
  or g27710 (n_14156, wc220, n_12072);
  not gc220 (wc220, \out_fifo[7][2] [0]);
  or g27711 (n_14115, wc221, n_12008);
  not gc221 (wc221, \out_fifo[2][1] [0]);
  or g27712 (n_14114, wc222, n_12007);
  not gc222 (wc222, \out_fifo[1][1] [0]);
  or g27713 (n_14112, wc223, n_12005);
  not gc223 (wc223, \out_fifo[3][1] [0]);
  or g27715 (n_14110, wc224, n_12070);
  not gc224 (wc224, \out_fifo[5][1] [0]);
  or g27716 (n_14109, wc225, n_12071);
  not gc225 (wc225, \out_fifo[6][1] [0]);
  or g27717 (n_14108, wc226, n_12072);
  not gc226 (wc226, \out_fifo[7][1] [0]);
  or g27718 (n_14067, wc227, n_12008);
  not gc227 (wc227, \out_fifo[2][0] [1]);
  nand g27719 (n_12034, n_11509, n_11511);
  or g27720 (n_14066, wc228, n_12007);
  not gc228 (wc228, \out_fifo[1][0] [1]);
  or g27721 (n_14064, wc229, n_12005);
  not gc229 (wc229, \out_fifo[3][0] [1]);
  or g27722 (n_14062, wc230, n_12070);
  not gc230 (wc230, \out_fifo[5][0] [1]);
  or g27723 (n_14061, wc231, n_12071);
  not gc231 (wc231, \out_fifo[6][0] [1]);
  or g27724 (n_14060, wc232, n_12072);
  not gc232 (wc232, \out_fifo[7][0] [1]);
  or g27725 (n_14019, wc233, n_12008);
  not gc233 (wc233, \out_fifo[2][0] [2]);
  or g27726 (n_14018, wc234, n_12007);
  not gc234 (wc234, \out_fifo[1][0] [2]);
  or g27727 (n_14016, wc235, n_12005);
  not gc235 (wc235, \out_fifo[3][0] [2]);
  or g27728 (n_14014, wc236, n_12070);
  not gc236 (wc236, \out_fifo[5][0] [2]);
  or g27729 (n_14013, wc237, n_12071);
  not gc237 (wc237, \out_fifo[6][0] [2]);
  or g27730 (n_14012, wc238, n_12072);
  not gc238 (wc238, \out_fifo[7][0] [2]);
  or g27731 (n_13971, wc239, n_12008);
  not gc239 (wc239, \out_fifo[2][0] [3]);
  or g27732 (n_13970, wc240, n_12007);
  not gc240 (wc240, \out_fifo[1][0] [3]);
  or g27733 (n_13968, wc241, n_12005);
  not gc241 (wc241, \out_fifo[3][0] [3]);
  or g27734 (n_13966, wc242, n_12070);
  not gc242 (wc242, \out_fifo[5][0] [3]);
  or g27735 (n_13965, wc243, n_12071);
  not gc243 (wc243, \out_fifo[6][0] [3]);
  or g27736 (n_13964, wc244, n_12072);
  not gc244 (wc244, \out_fifo[7][0] [3]);
  or g27737 (n_13923, wc245, n_12008);
  not gc245 (wc245, \out_fifo[2][0] [4]);
  or g27738 (n_13922, wc246, n_12007);
  not gc246 (wc246, \out_fifo[1][0] [4]);
  or g27739 (n_13920, wc247, n_12005);
  not gc247 (wc247, \out_fifo[3][0] [4]);
  or g27740 (n_13918, wc248, n_12070);
  not gc248 (wc248, \out_fifo[5][0] [4]);
  or g27741 (n_13917, wc249, n_12071);
  not gc249 (wc249, \out_fifo[6][0] [4]);
  or g27742 (n_13916, wc250, n_12072);
  not gc250 (wc250, \out_fifo[7][0] [4]);
  or g27743 (n_13875, wc251, n_12008);
  not gc251 (wc251, \out_fifo[2][0] [7]);
  or g27744 (n_13874, wc252, n_12007);
  not gc252 (wc252, \out_fifo[1][0] [7]);
  or g27745 (n_13872, wc253, n_12005);
  not gc253 (wc253, \out_fifo[3][0] [7]);
  or g27746 (n_13870, wc254, n_12070);
  not gc254 (wc254, \out_fifo[5][0] [7]);
  or g27747 (n_13869, wc255, n_12071);
  not gc255 (wc255, \out_fifo[6][0] [7]);
  or g27748 (n_13868, wc256, n_12072);
  not gc256 (wc256, \out_fifo[7][0] [7]);
  or g27749 (n_13395, wc257, n_11486);
  not gc257 (wc257, sh_reg_in[6]);
  or g27750 (n_13826, wc258, n_12007);
  not gc258 (wc258, \out_fifo[1][0] [5]);
  or g27751 (n_13824, wc259, n_12005);
  not gc259 (wc259, \out_fifo[3][0] [5]);
  or g27752 (n_13822, wc260, n_12070);
  not gc260 (wc260, \out_fifo[5][0] [5]);
  or g27753 (n_13821, wc261, n_12071);
  not gc261 (wc261, \out_fifo[6][0] [5]);
  or g27754 (n_13820, wc262, n_12072);
  not gc262 (wc262, \out_fifo[7][0] [5]);
  or g27755 (n_13779, wc263, n_12008);
  not gc263 (wc263, \out_fifo[2][0] [6]);
  or g27756 (n_13778, wc264, n_12007);
  not gc264 (wc264, \out_fifo[1][0] [6]);
  or g27757 (n_13776, wc265, n_12005);
  not gc265 (wc265, \out_fifo[3][0] [6]);
  or g27758 (n_13774, wc266, n_12070);
  not gc266 (wc266, \out_fifo[5][0] [6]);
  or g27759 (n_13773, wc267, n_12071);
  not gc267 (wc267, \out_fifo[6][0] [6]);
  or g27760 (n_13772, wc268, n_12072);
  not gc268 (wc268, \out_fifo[7][0] [6]);
  or g27761 (n_11564, data_stack_pointer[3], n_11563);
  or g27762 (n_13731, wc269, n_12008);
  not gc269 (wc269, \out_fifo[2][2] [8]);
  or g27763 (n_13730, wc270, n_12007);
  not gc270 (wc270, \out_fifo[1][2] [8]);
  or g27764 (n_13728, wc271, n_12005);
  not gc271 (wc271, \out_fifo[3][2] [8]);
  or g27765 (n_13726, wc272, n_12070);
  not gc272 (wc272, \out_fifo[5][2] [8]);
  or g27766 (n_13725, wc273, n_12071);
  not gc273 (wc273, \out_fifo[6][2] [8]);
  nand g27767 (n_16326, n_12192, n_11528);
  or g27768 (n_16327, n_12192, n_11528);
  nand g27769 (n_11529, n_16326, n_16327);
  or g27770 (n_13724, wc274, n_12072);
  not gc274 (wc274, \out_fifo[7][2] [8]);
  or g27771 (n_13683, wc275, n_12008);
  not gc275 (wc275, \out_fifo[2][0] [8]);
  or g27772 (n_13682, wc276, n_12007);
  not gc276 (wc276, \out_fifo[1][0] [8]);
  or g27773 (n_13680, wc277, n_12005);
  not gc277 (wc277, \out_fifo[3][0] [8]);
  or g27774 (n_13678, wc278, n_12070);
  not gc278 (wc278, \out_fifo[5][0] [8]);
  or g27775 (n_13677, wc279, n_12071);
  not gc279 (wc279, \out_fifo[6][0] [8]);
  or g27776 (n_13676, wc280, n_12072);
  not gc280 (wc280, \out_fifo[7][0] [8]);
  or g27777 (n_14402, wc281, n_11568);
  not gc281 (wc281, \data_stack_mem[6] [1]);
  or g27778 (n_13635, wc282, n_12008);
  not gc282 (wc282, \out_fifo[2][1] [1]);
  or g27779 (n_13634, wc283, n_12007);
  not gc283 (wc283, \out_fifo[1][1] [1]);
  or g27780 (n_13632, wc284, n_12005);
  not gc284 (wc284, \out_fifo[3][1] [1]);
  or g27781 (n_13630, wc285, n_12070);
  not gc285 (wc285, \out_fifo[5][1] [1]);
  nand g27782 (n_14395, n_12225, n_14394);
  or g27783 (n_13629, wc286, n_12071);
  not gc286 (wc286, \out_fifo[6][1] [1]);
  or g27784 (n_13628, wc287, n_12072);
  not gc287 (wc287, \out_fifo[7][1] [1]);
  nand g27785 (n_15742, n_11608, n_12244);
  or g27786 (n_12748, wc288, n_11563);
  not gc288 (wc288, \data_stack_mem[7] [4]);
  or g27787 (n_15079, wc289, n_11511);
  not gc289 (wc289, \data_stack_mem[0] [4]);
  or g27788 (n_13587, wc290, n_12008);
  not gc290 (wc290, \out_fifo[2][2] [9]);
  or g27789 (n_13586, wc291, n_12007);
  not gc291 (wc291, \out_fifo[1][2] [9]);
  or g27790 (n_11572, n_11516, n_14329);
  or g27791 (n_13584, wc292, n_12005);
  not gc292 (wc292, \out_fifo[3][2] [9]);
  or g27792 (n_13582, wc293, n_12070);
  not gc293 (wc293, \out_fifo[5][2] [9]);
  or g27793 (n_13581, wc294, n_12071);
  not gc294 (wc294, \out_fifo[6][2] [9]);
  or g27794 (n_12751, wc295, n_11563);
  not gc295 (wc295, \data_stack_mem[7] [2]);
  or g27795 (n_13580, wc296, n_12072);
  not gc296 (wc296, \out_fifo[7][2] [9]);
  or g27796 (n_14854, wc297, n_11511);
  not gc297 (wc297, \data_stack_mem[0] [2]);
  or g27797 (n_13539, wc298, n_12008);
  not gc298 (wc298, \out_fifo[2][1] [2]);
  or g27798 (n_13538, wc299, n_12007);
  not gc299 (wc299, \out_fifo[1][1] [2]);
  or g27799 (n_12730, wc300, n_11563);
  not gc300 (wc300, \data_stack_mem[7] [7]);
  or g27800 (n_13536, wc301, n_12005);
  not gc301 (wc301, \out_fifo[3][1] [2]);
  or g27801 (n_15343, wc302, n_11511);
  not gc302 (wc302, \data_stack_mem[0] [7]);
  or g27802 (n_13534, wc303, n_12070);
  not gc303 (wc303, \out_fifo[5][1] [2]);
  or g27803 (n_13533, wc304, n_12071);
  not gc304 (wc304, \out_fifo[6][1] [2]);
  or g27804 (n_13532, wc305, n_12072);
  not gc305 (wc305, \out_fifo[7][1] [2]);
  or g27805 (n_13491, wc306, n_12008);
  not gc306 (wc306, \out_fifo[2][1] [3]);
  or g27806 (n_13359, wc307, n_11486);
  not gc307 (wc307, sh_reg_in[1]);
  nand g27807 (n_13360, \data_stack_mem[8] [1], n_11484);
  or g27808 (n_13365, wc308, n_11486);
  not gc308 (wc308, sh_reg_in[3]);
  nand g27809 (n_13366, \data_stack_mem[8] [3], n_11484);
  or g27810 (n_13371, wc309, n_11486);
  not gc309 (wc309, sh_reg_in[5]);
  nand g27811 (n_13372, \data_stack_mem[8] [5], n_11484);
  or g27812 (n_13377, wc310, n_11486);
  not gc310 (wc310, sh_reg_in[7]);
  nand g27813 (n_13378, \data_stack_mem[8] [7], n_11484);
  or g27814 (n_13383, wc311, n_11486);
  not gc311 (wc311, sh_reg_in[0]);
  nand g27815 (n_13384, \data_stack_mem[8] [0], n_11484);
  or g27816 (n_13389, wc312, n_11486);
  not gc312 (wc312, sh_reg_in[2]);
  nand g27817 (n_13390, \data_stack_mem[8] [2], n_11484);
  or g27818 (n_13490, wc313, n_12007);
  not gc313 (wc313, \out_fifo[1][1] [3]);
  or g27819 (n_14521, wc314, n_11511);
  not gc314 (wc314, \data_stack_mem[0] [0]);
  or g27820 (n_12006, out_fifo_read_pointer[0], n_13111);
  or g27821 (n_12742, wc315, n_11563);
  not gc315 (wc315, \data_stack_mem[7] [6]);
  or g27822 (n_13488, wc316, n_12005);
  not gc316 (wc316, \out_fifo[3][1] [3]);
  or g27823 (n_15259, wc317, n_11511);
  not gc317 (wc317, \data_stack_mem[0] [6]);
  or g27824 (n_13486, wc318, n_12070);
  not gc318 (wc318, \out_fifo[5][1] [3]);
  or g27825 (n_13485, wc319, n_12071);
  not gc319 (wc319, \out_fifo[6][1] [3]);
  or g27826 (n_13484, wc320, n_12072);
  not gc320 (wc320, \out_fifo[7][1] [3]);
  or g27827 (n_12073, out_fifo_read_pointer[0], n_13114);
  nand g27830 (n_14323, n_12244, n_14322);
  or g27833 (n_12757, wc321, n_11563);
  not gc321 (wc321, \data_stack_mem[7] [1]);
  or g27834 (n_13449, wc322, n_11896);
  not gc322 (wc322, sh_reg_in[7]);
  or g27835 (n_14728, wc323, n_11511);
  not gc323 (wc323, \data_stack_mem[0] [1]);
  or g27836 (n_13443, wc324, n_11896);
  not gc324 (wc324, sh_reg_in[6]);
  or g27837 (n_13437, wc325, n_11896);
  not gc325 (wc325, sh_reg_in[5]);
  or g27839 (n_13431, wc326, n_11896);
  not gc326 (wc326, sh_reg_in[4]);
  nand g27840 (n_15736, n_12278, n_11577);
  or g27841 (n_12745, wc327, n_11563);
  not gc327 (wc327, \data_stack_mem[7] [5]);
  or g27842 (n_15175, wc328, n_11511);
  not gc328 (wc328, \data_stack_mem[0] [5]);
  or g27843 (n_13425, wc329, n_11896);
  not gc329 (wc329, sh_reg_in[3]);
  or g27845 (n_13419, wc330, n_11896);
  not gc330 (wc330, sh_reg_in[2]);
  or g27846 (n_13413, wc331, n_11896);
  not gc331 (wc331, sh_reg_in[1]);
  or g27847 (n_12754, wc332, n_11563);
  not gc332 (wc332, \data_stack_mem[7] [3]);
  or g27848 (n_14932, wc333, n_11511);
  not gc333 (wc333, \data_stack_mem[0] [3]);
  or g27850 (n_13407, wc334, n_11896);
  not gc334 (wc334, sh_reg_in[0]);
  nand g27851 (n_13402, \data_stack_mem[8] [4], n_11484);
  or g27852 (n_13401, wc335, n_11486);
  not gc335 (wc335, sh_reg_in[4]);
  nand g27853 (n_13396, \data_stack_mem[8] [6], n_11484);
  or g27854 (n_13827, wc336, n_12008);
  not gc336 (wc336, \out_fifo[2][0] [5]);
  nand g27855 (n_15666, \out_fifo[7][1] [3], n_11498);
  nand g27856 (n_15672, \out_fifo[3][1] [3], n_11543);
  nand g27857 (n_15678, \out_fifo[7][1] [0], n_11498);
  nand g27858 (n_14964, \out_fifo[4][0] [4], n_11556);
  nand g27859 (n_13026, \out_fifo[3][2] [0], n_11543);
  or g27860 (n_11896, data_stack_pointer[3], n_12874);
  nand g27861 (n_14971, \out_fifo[5][0] [4], n_11560);
  nand g27862 (n_12023, n_11544, n_13039);
  nand g27863 (n_13044, n_11552, \out_fifo[2][2] [1]);
  nand g27864 (n_15684, \out_fifo[0][1] [0], n_11535);
  nand g27865 (n_15661, \out_fifo[5][1] [3], n_11560);
  nand g27866 (n_15690, \out_fifo[6][1] [0], n_11540);
  nand g27867 (n_15696, \out_fifo[1][1] [0], n_11548);
  or g27868 (n_11655, n_11654, n_12715);
  nand g27869 (n_15654, \out_fifo[4][1] [3], n_11556);
  nand g27870 (n_12823, n_12215, n_12822);
  nand g27871 (n_15642, \out_fifo[1][1] [3], n_11548);
  nand g27872 (n_14982, \out_fifo[7][0] [4], n_11498);
  or g27873 (n_13045, n_11538, n_12028);
  nand g27874 (n_15636, \out_fifo[6][1] [3], n_11540);
  nand g27875 (n_13050, n_11560, \out_fifo[5][2] [1]);
  nand g27876 (n_15630, \out_fifo[0][1] [3], n_11535);
  nand g27877 (n_15615, \out_fifo[3][0] [0], n_11543);
  nand g27878 (n_15609, \out_fifo[3][1] [2], n_11543);
  or g27879 (n_13051, n_11546, n_11908);
  nand g27881 (n_13056, n_11535, \out_fifo[0][2] [1]);
  or g27883 (n_13057, n_11532, n_12028);
  nand g27884 (n_13062, n_11543, \out_fifo[3][2] [1]);
  nand g27885 (n_15702, \out_fifo[2][1] [0], n_11552);
  nand g27886 (n_15604, \out_fifo[5][0] [0], n_11560);
  or g27887 (n_13063, n_11495, n_12028);
  nand g27888 (n_13068, n_11548, \out_fifo[1][2] [1]);
  or g27889 (n_13069, n_11546, n_12028);
  nand g27890 (n_15597, \out_fifo[4][0] [0], n_11556);
  nand g27891 (n_15591, \out_fifo[2][0] [0], n_11552);
  nand g27892 (n_15585, \out_fifo[1][0] [0], n_11548);
  nand g27893 (n_13074, n_11498, \out_fifo[7][2] [1]);
  nand g27894 (n_15579, \out_fifo[6][0] [0], n_11540);
  nand g27895 (n_15573, \out_fifo[0][0] [0], n_11535);
  nand g27896 (n_15567, \out_fifo[7][0] [0], n_11498);
  nand g27897 (n_15561, \out_fifo[7][1] [2], n_11498);
  nand g27898 (n_14988, \out_fifo[3][0] [4], n_11543);
  or g27899 (n_13075, n_11495, n_11908);
  nand g27900 (n_13080, n_11540, \out_fifo[6][2] [1]);
  or g27901 (n_13081, n_11538, n_11908);
  or g27902 (n_11912, n_11871, n_11507);
  nand g27903 (n_13086, n_11556, \out_fifo[4][2] [1]);
  or g27904 (n_13087, n_11532, n_11908);
  nand g27905 (n_15087, \out_fifo[0][0] [5], n_11535);
  nand g27906 (n_11484, n_12117, n_13099);
  or g27907 (n_13317, wc337, n_11992);
  not gc337 (wc337, sh_reg_in[1]);
  nand g27908 (n_13105, n_13104, n_12117);
  nand g27909 (n_11952, n_12654, n_12655);
  or g27910 (n_11980, n_11871, n_11968);
  nand g27911 (n_13108, n_12333, rst_n);
  or g27912 (n_13119, wc338, n_11867);
  not gc338 (wc338, sh_reg_in[7]);
  nand g27913 (n_15556, \out_fifo[5][1] [2], n_11560);
  nand g27914 (n_15549, \out_fifo[4][1] [2], n_11556);
  or g27915 (n_13125, wc339, n_11867);
  not gc339 (wc339, sh_reg_in[4]);
  or g27916 (n_13131, wc340, n_11867);
  not gc340 (wc340, sh_reg_in[0]);
  or g27917 (n_13137, wc341, n_11867);
  not gc341 (wc341, sh_reg_in[5]);
  or g27918 (n_13143, wc342, n_11867);
  not gc342 (wc342, sh_reg_in[1]);
  nand g27919 (n_14322, \data_stack_mem[2] [2], n_11604);
  nand g27921 (n_15708, \out_fifo[4][1] [0], n_11556);
  nand g27922 (n_15715, \out_fifo[5][1] [0], n_11560);
  or g27923 (n_13114, out_fifo_read_pointer[1], n_12003);
  nand g27924 (n_15720, \out_fifo[3][1] [0], n_11543);
  or g27925 (n_13149, wc343, n_11867);
  not gc343 (wc343, sh_reg_in[2]);
  nand g27926 (n_12305, n_12840, n_12841);
  nand g27927 (n_15648, \out_fifo[2][1] [3], n_11552);
  or g27928 (n_14334, wc344, n_11969);
  not gc344 (wc344, sh_reg_in[1]);
  or g27929 (n_13155, wc345, n_11867);
  not gc345 (wc345, sh_reg_in[3]);
  nand g27930 (n_12027, n_12681, n_12682);
  or g27931 (n_14340, wc346, n_11969);
  not gc346 (wc346, sh_reg_in[7]);
  or g27932 (n_13161, wc347, n_11867);
  not gc347 (wc347, sh_reg_in[6]);
  or g27933 (n_14346, wc348, n_11969);
  not gc348 (wc348, sh_reg_in[4]);
  or g27934 (n_13168, wc349, n_11883);
  not gc349 (wc349, sh_reg_in[7]);
  or g27935 (n_13174, wc350, n_11883);
  not gc350 (wc350, sh_reg_in[6]);
  or g27936 (n_13180, wc351, n_11883);
  not gc351 (wc351, sh_reg_in[5]);
  or g27937 (n_13186, wc352, n_11883);
  not gc352 (wc352, sh_reg_in[4]);
  nand g27938 (n_15543, \out_fifo[2][1] [2], n_11552);
  nand g27939 (n_15733, \data_stack_mem[0] [3], n_12215);
  nand g27940 (n_15537, \out_fifo[1][1] [2], n_11548);
  nand g27941 (n_15531, \out_fifo[6][1] [2], n_11540);
  nand g27942 (n_15525, \out_fifo[0][1] [2], n_11535);
  nand g27943 (n_15510, \out_fifo[3][1] [1], n_11543);
  nand g27944 (n_15504, \out_fifo[7][1] [1], n_11498);
  nand g27945 (n_15498, \out_fifo[3][1] [4], n_11543);
  nand g27946 (n_15492, \out_fifo[7][1] [4], n_11498);
  or g27947 (n_13111, out_fifo_read_pointer[1], n_12004);
  or g27948 (n_14352, wc353, n_11969);
  not gc353 (wc353, sh_reg_in[6]);
  nand g27949 (n_11954, n_12762, n_12763);
  or g27950 (n_12005, n_12001, n_12004);
  or g27951 (n_12007, n_12004, n_11861);
  or g27952 (n_12008, n_12004, n_11862);
  or g27953 (n_13353, wc354, n_11992);
  not gc354 (wc354, sh_reg_in[2]);
  or g27954 (n_11522, n_12865, n_11510);
  or g27955 (n_13192, wc355, n_11883);
  not gc355 (wc355, sh_reg_in[3]);
  nand g27956 (n_15487, \out_fifo[5][1] [4], n_11560);
  nand g27957 (n_15480, \out_fifo[4][1] [4], n_11556);
  nand g27958 (n_15474, \out_fifo[2][1] [4], n_11552);
  nand g27959 (n_15468, \out_fifo[1][1] [4], n_11548);
  or g27960 (n_14358, wc356, n_11969);
  not gc356 (wc356, sh_reg_in[5]);
  nand g27961 (n_15462, \out_fifo[6][1] [4], n_11540);
  nand g27962 (n_15456, \out_fifo[0][1] [4], n_11535);
  nand g27963 (n_15451, \out_fifo[5][1] [1], n_11560);
  or g27964 (n_13198, wc357, n_11883);
  not gc357 (wc357, sh_reg_in[2]);
  nand g27965 (n_15444, \out_fifo[4][1] [1], n_11556);
  nand g27966 (n_15438, \out_fifo[2][1] [1], n_11552);
  nand g27967 (n_15432, \out_fifo[1][1] [1], n_11548);
  nand g27968 (n_15426, \out_fifo[6][1] [1], n_11540);
  nand g27969 (n_15420, \out_fifo[0][1] [1], n_11535);
  nand g27970 (n_15393, \out_fifo[3][0] [8], n_11543);
  nand g27971 (n_15387, \out_fifo[7][0] [8], n_11498);
  or g27972 (n_13347, wc358, n_11992);
  not gc358 (wc358, sh_reg_in[3]);
  nand g27973 (n_12365, n_11505, n_12616);
  or g27974 (n_14364, wc359, n_11969);
  not gc359 (wc359, sh_reg_in[2]);
  or g27975 (n_13341, wc360, n_11992);
  not gc360 (wc360, sh_reg_in[4]);
  or g27976 (n_13335, wc361, n_11992);
  not gc361 (wc361, sh_reg_in[0]);
  or g27977 (n_13329, wc362, n_11992);
  not gc362 (wc362, sh_reg_in[6]);
  or g27978 (n_13323, wc363, n_11992);
  not gc363 (wc363, sh_reg_in[5]);
  or g27979 (n_12070, n_11861, n_12003);
  or g27980 (n_12071, n_11862, n_12003);
  or g27981 (n_13204, wc364, n_11883);
  not gc364 (wc364, sh_reg_in[1]);
  or g27982 (n_12072, n_12001, n_12003);
  or g27983 (n_14370, wc365, n_11969);
  not gc365 (wc365, sh_reg_in[0]);
  or g27984 (n_13210, wc366, n_11883);
  not gc366 (wc366, sh_reg_in[0]);
  or g27985 (n_14376, wc367, n_11969);
  not gc367 (wc367, sh_reg_in[3]);
  nand g27986 (n_15382, \out_fifo[5][0] [8], n_11560);
  nand g27987 (n_15375, \out_fifo[4][0] [8], n_11556);
  nand g27988 (n_15369, \out_fifo[2][0] [8], n_11552);
  nand g27989 (n_15363, \out_fifo[1][0] [8], n_11548);
  nand g27990 (n_15357, \out_fifo[6][0] [8], n_11540);
  nand g27991 (n_15351, \out_fifo[0][0] [8], n_11535);
  nand g27992 (n_15309, \out_fifo[3][0] [7], n_11543);
  or g27993 (n_13311, wc368, n_11992);
  not gc368 (wc368, sh_reg_in[7]);
  nand g27994 (n_16328, n_12280, n_11576);
  or g27995 (n_16329, n_12280, n_11576);
  nand g27996 (n_11577, n_16328, n_16329);
  nand g27997 (n_15303, \out_fifo[7][0] [7], n_11498);
  nand g27998 (n_15298, \out_fifo[5][0] [7], n_11560);
  nand g27999 (n_15291, \out_fifo[4][0] [7], n_11556);
  nand g28000 (n_14526, \out_fifo[0][0] [1], n_11535);
  nand g28001 (n_14532, \out_fifo[6][0] [1], n_11540);
  nand g28002 (n_11884, n_12117, n_11485);
  nand g28003 (n_14538, \out_fifo[1][0] [1], n_11548);
  nand g28004 (n_14544, \out_fifo[2][0] [1], n_11552);
  nand g28005 (n_14550, \out_fifo[4][0] [1], n_11556);
  nand g28006 (n_14557, \out_fifo[5][0] [1], n_11560);
  nand g28007 (n_15285, \out_fifo[2][0] [7], n_11552);
  nand g28008 (n_14568, \out_fifo[7][0] [1], n_11498);
  nand g28009 (n_14574, \out_fifo[3][0] [1], n_11543);
  nand g28010 (n_14736, \out_fifo[0][0] [2], n_11535);
  nand g28011 (n_15279, \out_fifo[1][0] [7], n_11548);
  nand g28012 (n_14742, \out_fifo[6][0] [2], n_11540);
  nand g28013 (n_15273, \out_fifo[6][0] [7], n_11540);
  nand g28014 (n_14748, \out_fifo[1][0] [2], n_11548);
  nand g28015 (n_15267, \out_fifo[0][0] [7], n_11535);
  nand g28016 (n_15225, \out_fifo[3][0] [6], n_11543);
  nand g28017 (n_15219, \out_fifo[7][0] [6], n_11498);
  nand g28018 (n_15214, \out_fifo[5][0] [6], n_11560);
  nand g28019 (n_15207, \out_fifo[4][0] [6], n_11556);
  nand g28020 (n_15201, \out_fifo[2][0] [6], n_11552);
  nand g28021 (n_15195, \out_fifo[1][0] [6], n_11548);
  nand g28022 (n_14754, \out_fifo[2][0] [2], n_11552);
  nand g28023 (n_14760, \out_fifo[4][0] [2], n_11556);
  nand g28024 (n_14767, \out_fifo[5][0] [2], n_11560);
  nand g28025 (n_14784, \out_fifo[7][0] [2], n_11498);
  nand g28026 (n_14790, \out_fifo[3][0] [2], n_11543);
  nand g28027 (n_14329, n_12238, n_14328);
  nand g28028 (n_14862, \out_fifo[0][0] [3], n_11535);
  nand g28029 (n_14868, \out_fifo[6][0] [3], n_11540);
  nand g28031 (n_14874, \out_fifo[1][0] [3], n_11548);
  nand g28032 (n_15189, \out_fifo[6][0] [6], n_11540);
  nand g28033 (n_14880, \out_fifo[2][0] [3], n_11552);
  nand g28034 (n_14886, \out_fifo[4][0] [3], n_11556);
  nand g28036 (n_15183, \out_fifo[0][0] [6], n_11535);
  nand g28037 (n_15129, \out_fifo[3][0] [5], n_11543);
  nand g28038 (n_15123, \out_fifo[7][0] [5], n_11498);
  nand g28039 (n_14893, \out_fifo[5][0] [3], n_11560);
  nand g28040 (n_15118, \out_fifo[5][0] [5], n_11560);
  nand g28041 (n_14910, \out_fifo[7][0] [3], n_11498);
  nand g28042 (n_15111, \out_fifo[4][0] [5], n_11556);
  nand g28043 (n_15105, \out_fifo[2][0] [5], n_11552);
  nand g28044 (n_14916, \out_fifo[3][0] [3], n_11543);
  nand g28045 (n_12883, n_12881, n_12882);
  nand g28046 (n_15099, \out_fifo[1][0] [5], n_11548);
  nand g28047 (n_12888, \out_fifo[0][2] [0], n_11535);
  nand g28048 (n_12894, \out_fifo[6][2] [0], n_11540);
  nand g28049 (n_12900, \out_fifo[1][2] [0], n_11548);
  nand g28050 (n_14940, \out_fifo[0][0] [4], n_11535);
  nand g28051 (n_12906, \out_fifo[2][2] [0], n_11552);
  nand g28052 (n_12912, \out_fifo[4][2] [0], n_11556);
  nand g28053 (n_12919, \out_fifo[5][2] [0], n_11560);
  or g28054 (n_14394, wc369, n_11569);
  not gc369 (wc369, \data_stack_mem[5] [1]);
  nand g28055 (n_14946, \out_fifo[6][0] [4], n_11540);
  or g28056 (n_12924, wc370, n_12044);
  not gc370 (wc370, sh_reg_in[7]);
  or g28057 (n_12930, wc371, n_12044);
  not gc371 (wc371, sh_reg_in[5]);
  or g28058 (n_12936, wc372, n_12044);
  not gc372 (wc372, sh_reg_in[6]);
  or g28059 (n_12942, wc373, n_12044);
  not gc373 (wc373, sh_reg_in[3]);
  or g28060 (n_12948, wc374, n_12044);
  not gc374 (wc374, sh_reg_in[4]);
  or g28061 (n_12954, wc375, n_12044);
  not gc375 (wc375, sh_reg_in[2]);
  or g28062 (n_12960, wc376, n_12044);
  not gc376 (wc376, sh_reg_in[1]);
  or g28063 (n_12966, wc377, n_12044);
  not gc377 (wc377, sh_reg_in[0]);
  nand g28064 (n_12972, \out_fifo[7][2] [8], n_11498);
  nand g28065 (n_12978, \out_fifo[3][2] [8], n_11543);
  nand g28066 (n_14952, \out_fifo[1][0] [4], n_11548);
  nand g28067 (n_15093, \out_fifo[6][0] [5], n_11540);
  nand g28068 (n_12984, \out_fifo[7][2] [0], n_11498);
  nand g28069 (n_12990, \out_fifo[0][2] [8], n_11535);
  nand g28070 (n_12996, \out_fifo[6][2] [8], n_11540);
  nand g28071 (n_13002, \out_fifo[1][2] [8], n_11548);
  nand g28072 (n_13008, \out_fifo[2][2] [8], n_11552);
  nand g28073 (n_13014, \out_fifo[4][2] [8], n_11556);
  nand g28074 (n_16330, n_12197, n_11527);
  or g28075 (n_16331, n_12197, n_11527);
  nand g28076 (n_11528, n_16330, n_16331);
  nand g28077 (n_13021, \out_fifo[5][2] [8], n_11560);
  nand g28078 (n_14958, \out_fifo[2][0] [4], n_11552);
  or g28079 (n_11969, n_12805, n_11881);
  or g28081 (n_11479, n_11478, wc378);
  not gc378 (wc378, n_12814);
  or g28082 (n_11867, n_11866, n_11507);
  nand g28083 (n_11543, n_11496, n_12029);
  or g28086 (n_12637, wc379, n_11510);
  not gc379 (wc379, n_12367);
  or g28087 (n_11536, n_11534, wc380);
  not gc380 (wc380, rst_n);
  or g28088 (n_12655, n_12653, wc381);
  not gc381 (wc381, rst_n);
  nand g28089 (n_12640, n_11502, n_11510);
  nand g28090 (n_11869, n_12786, n_12787);
  or g28091 (n_11871, data_stack_pointer[0], n_11868);
  or g28092 (n_12333, wc382, n_11970);
  not gc382 (wc382, n_11507);
  or g28093 (n_11883, n_11483, n_11882);
  nand g28094 (n_11498, n_11496, n_11907);
  or g28095 (n_11688, n_11687, n_12775);
  or g28096 (n_11506, n_11502, n_11504);
  nand g28097 (n_12025, n_12672, n_12673);
  or g28098 (n_11557, n_11555, wc383);
  not gc383 (wc383, rst_n);
  or g28099 (n_12044, n_12805, n_11485);
  or g28100 (n_11505, wc384, n_11502);
  not gc384 (wc384, n_11504);
  or g28101 (n_14328, wc385, n_11571);
  not gc385 (wc385, \data_stack_mem[4] [1]);
  or g28103 (n_11587, n_11586, n_12772);
  nand g28104 (n_12822, \data_stack_mem[1] [3], n_11643);
  nand g28105 (n_12881, n_11970, rst_n);
  nand g28106 (n_11604, n_12737, n_15730);
  or g28107 (n_12874, n_11483, n_11485);
  or g28109 (n_11966, n_11478, wc386);
  not gc386 (wc386, n_12859);
  or g28110 (n_11967, n_11478, wc387);
  not gc387 (wc387, n_12856);
  or g28111 (n_11965, n_11478, wc388);
  not gc388 (wc388, n_12853);
  nand g28112 (n_11556, n_12850, n_11907);
  nand g28113 (n_11535, n_12029, n_12850);
  nand g28114 (n_16332, n_12231, n_11526);
  or g28115 (n_16333, n_12231, n_11526);
  nand g28116 (n_11527, n_16332, n_16333);
  nand g28117 (n_12762, n_12354, rst_n);
  nand g28118 (n_11953, n_12726, n_12727);
  nand g28119 (n_16334, n_11607, \data_stack_mem[0] [2]);
  or g28120 (n_16335, n_11607, \data_stack_mem[0] [2]);
  nand g28121 (n_11608, n_16334, n_16335);
  or g28122 (n_11541, n_11539, wc389);
  not gc389 (wc389, rst_n);
  nand g28123 (n_12003, out_fifo_read_pointer[2], n_11478);
  or g28124 (n_12004, out_fifo_read_pointer[2], wc390);
  not gc390 (wc390, n_11478);
  or g28125 (n_12865, n_11521, n_12864);
  or g28126 (n_11549, n_11547, wc391);
  not gc391 (wc391, rst_n);
  nand g28127 (n_11548, n_12847, n_12029);
  or g28128 (n_12616, \data_stack_mem[8] [0], n_11502);
  nand g28129 (n_11560, n_11907, n_12847);
  or g28130 (n_11561, n_11559, wc392);
  not gc392 (wc392, rst_n);
  nand g28131 (n_11540, n_12844, n_11907);
  nand g28132 (n_11552, n_12029, n_12844);
  or g28133 (n_12280, n_12739, wc393);
  not gc393 (wc393, n_11517);
  nand g28134 (n_12117, rst_n, n_11483);
  nand g28135 (n_12024, n_12549, n_12550);
  or g28136 (n_11553, n_11551, wc394);
  not gc394 (wc394, rst_n);
  or g28138 (n_12682, n_12680, wc395);
  not gc395 (wc395, rst_n);
  or g28139 (n_12028, out_fifo_write_pointer[2], n_12118);
  or g28140 (n_11992, n_11866, n_11968);
  or g28142 (n_12654, data_stack_pointer[2], n_12652);
  or g28143 (n_11480, n_11478, wc396);
  not gc396 (wc396, n_12817);
  or g28144 (n_11544, n_11894, wc397);
  not gc397 (wc397, rst_n);
  or g28145 (n_11500, n_11893, wc398);
  not gc398 (wc398, rst_n);
  or g28146 (n_11866, n_11512, n_11865);
  or g28147 (n_11868, wc399, n_11865);
  not gc399 (wc399, data_stack_pointer[1]);
  or g28150 (n_13039, wc400, n_12114);
  not gc400 (wc400, n_12337);
  or g28151 (n_11893, n_11495, n_11497);
  not g28152 (n_16336, n_11893);
  or g28153 (n_11722, n_11721, n_12778);
  or g28154 (n_12831, wc401, n_11573);
  not gc401 (wc401, \data_stack_mem[3] [1]);
  or g28155 (n_11894, n_11495, n_11533);
  not g28156 (n_16337, n_11894);
  nand g28157 (n_15730, n_12295, n_11576);
  or g28158 (n_11586, n_12694, wc402);
  not gc402 (wc402, n_12138);
  nand g28159 (n_12839, n_11573, \data_stack_mem[3] [1]);
  nand g28160 (n_11478, n_12798, n_12799);
  or g28161 (n_11756, n_11755, n_12769);
  or g28162 (n_11607, n_12661, wc403);
  not gc403 (wc403, n_11508);
  or g28163 (n_11521, n_11520, n_12766);
  or g28164 (n_12840, n_11573, n_12138);
  or g28165 (n_11510, sh_reg_in[4], n_12490);
  or g28166 (n_12118, n_11509, n_12718);
  nand g28167 (n_12739, n_12295, n_12737);
  nand g28170 (n_12029, n_11533, rst_n);
  or g28172 (n_11687, n_12697, wc404);
  not gc404 (wc404, n_12152);
  nand g28173 (n_11907, n_11497, rst_n);
  or g28174 (n_12805, n_11482, n_11968);
  or g28175 (n_12763, wc405, n_11906);
  not gc405 (wc405, out_fifo_write_pointer[1]);
  or g28176 (n_12727, wc406, n_11906);
  not gc406 (wc406, out_fifo_write_pointer[0]);
  or g28177 (n_12726, n_12725, wc407);
  not gc407 (wc407, rst_n);
  nand g28178 (n_12520, n_12517, n_12518);
  nand g28179 (n_12680, n_11951, data_stack_pointer[3]);
  or g28180 (n_12681, wc408, n_12175);
  not gc408 (wc408, n_12356);
  nand g28181 (n_11470, n_12525, n_12526);
  or g28182 (n_12672, wc409, n_12175);
  not gc409 (wc409, n_12355);
  or g28183 (n_12550, n_12548, wc410);
  not gc410 (wc410, rst_n);
  nand g28184 (n_12354, n_11538, n_12664);
  or g28185 (n_12549, out_fifo_read_pointer[2], n_12547);
  or g28186 (n_12652, n_11512, n_12651);
  nand g28187 (n_12026, n_12582, n_12583);
  nand g28188 (n_12653, n_11951, data_stack_pointer[2]);
  nand g28189 (n_16338, n_12262, n_11525);
  or g28190 (n_16339, n_12262, n_11525);
  nand g28191 (n_11526, n_16338, n_16339);
  nand g28192 (n_11643, n_12660, n_15727);
  or g28194 (n_13775, wc411, n_11457);
  not gc411 (wc411, sh_reg_out[5]);
  nand g28195 (n_11948, n_12612, n_12613);
  nand g28196 (n_12356, n_12600, n_12601);
  or g28197 (n_11951, n_11481, wc412);
  not gc412 (wc412, n_12634);
  or g28198 (n_12651, n_11864, n_11950);
  nand g28199 (n_16340, n_12261, n_11524);
  or g28200 (n_16341, n_12261, n_11524);
  nand g28201 (n_11525, n_16340, n_16341);
  nand g28202 (n_12355, n_12591, n_12592);
  or g28205 (n_13823, wc413, n_11457);
  not gc413 (wc413, sh_reg_out[4]);
  or g28208 (n_12582, n_11481, n_12581);
  or g28209 (n_13727, wc414, n_11457);
  not gc414 (wc414, sh_reg_out[27]);
  or g28210 (n_12664, n_11546, n_11905);
  or g28213 (n_12547, n_12001, n_12113);
  nand g28214 (n_15727, \data_stack_mem[0] [2], n_12213);
  or g28215 (n_12673, n_12671, wc415);
  not gc415 (wc415, rst_n);
  nand g28216 (n_12548, n_12362, out_fifo_read_pointer[2]);
  or g28217 (n_13871, wc416, n_11457);
  not gc416 (wc416, sh_reg_out[6]);
  or g28218 (n_13679, wc417, n_11457);
  not gc417 (wc417, sh_reg_out[7]);
  or g28219 (n_12525, out_fifo_read_pointer[0], n_12113);
  or g28220 (n_12518, wc418, n_12112);
  not gc418 (wc418, out_fifo_read_pointer[1]);
  or g28221 (n_12517, n_11861, n_12113);
  or g28222 (n_12725, n_11905, out_fifo_write_pointer[0]);
  or g28223 (n_11477, n_12508, wc419);
  not gc419 (wc419, rst_n);
  or g28226 (n_13631, wc420, n_11457);
  not gc420 (wc420, sh_reg_out[10]);
  or g28227 (n_13919, wc421, n_11457);
  not gc421 (wc421, sh_reg_out[3]);
  or g28238 (n_12697, wc422, n_11686);
  not gc422 (wc422, n_12387);
  or g28239 (n_12337, n_11495, n_11905);
  or g28242 (n_12814, wc423, n_11457);
  not gc423 (wc423, dout_valid);
  or g28243 (n_13967, wc424, n_11457);
  not gc424 (wc424, sh_reg_out[2]);
  or g28244 (n_12493, sh_reg_in[0], n_11501);
  or g28245 (n_12737, wc425, n_11574);
  not gc425 (wc425, \data_stack_mem[2] [1]);
  or g28246 (n_12817, sh_reg_out_bit_counter[0], n_11457);
  or g28247 (n_13583, wc426, n_11457);
  not gc426 (wc426, sh_reg_out[28]);
  or g28248 (n_12711, n_11619, n_12710);
  or g28250 (n_11813, n_11812, n_12703);
  or g28253 (n_13535, wc427, n_11457);
  not gc427 (wc427, sh_reg_out[11]);
  or g28254 (n_11520, n_11519, n_12688);
  or g28255 (n_14015, wc428, n_11457);
  not gc428 (wc428, sh_reg_out[1]);
  or g28256 (n_11755, n_11754, n_12691);
  or g28257 (n_12799, out_fifo_read_pointer[2], n_12797);
  nand g28259 (n_12661, n_12213, n_12660);
  or g28264 (n_13487, wc429, n_11457);
  not gc429 (wc429, sh_reg_out[12]);
  or g28265 (n_12798, wc430, n_12172);
  not gc430 (wc430, n_12329);
  or g28266 (n_14063, wc431, n_11457);
  not gc431 (wc431, sh_reg_out[0]);
  or g28269 (n_12694, wc432, n_11585);
  not gc432 (wc432, n_12382);
  or g28270 (n_14111, wc433, n_11457);
  not gc433 (wc433, sh_reg_out[9]);
  or g28271 (n_14159, wc434, n_11457);
  not gc434 (wc434, sh_reg_out[19]);
  nand g28272 (n_11906, rst_n, n_11905);
  or g28273 (n_11721, n_11720, n_12700);
  or g28274 (n_14207, wc435, n_11457);
  not gc435 (wc435, sh_reg_out[13]);
  or g28275 (n_14255, wc436, n_11457);
  not gc436 (wc436, sh_reg_out[20]);
  nand g28276 (n_12787, n_12253, rst_n);
  or g28277 (n_12630, n_12629, wc437);
  not gc437 (wc437, n_12148);
  or g28278 (n_11865, sh_reg_in[8], n_11864);
  or g28279 (n_12526, wc438, n_12112);
  not gc438 (wc438, out_fifo_read_pointer[0]);
  or g28280 (n_11501, sh_reg_in[6], n_12460);
  nand g28281 (n_12778, n_12397, n_12396);
  nand g28282 (n_11949, n_12558, n_12559);
  nand g28283 (n_12864, n_12375, n_12374);
  or g28284 (n_12581, n_11950, n_11485);
  nand g28286 (n_12629, n_12409, n_12408);
  nand g28287 (n_11754, n_12381, n_12380);
  nand g28288 (n_16355, n_11575, \data_stack_mem[0] [1]);
  or g28289 (n_16356, n_11575, \data_stack_mem[0] [1]);
  nand g28290 (n_11576, n_16355, n_16356);
  or g28291 (n_12591, n_11481, n_12590);
  nand g28292 (n_11686, n_12391, n_12390);
  nand g28293 (n_12691, n_12379, n_12378);
  nand g28294 (n_11457, n_11456, rst_n);
  nand g28295 (n_12715, n_12407, n_12406);
  nand g28296 (n_12775, n_12395, n_12394);
  nand g28297 (n_12769, n_12377, n_12376);
  nand g28298 (n_12660, \data_stack_mem[1] [2], n_11606);
  nand g28299 (n_12508, n_11481, n_12507);
  nand g28301 (n_16357, n_12266, n_11523);
  or g28302 (n_16358, n_12266, n_11523);
  nand g28303 (n_11524, n_16357, n_16358);
  or g28304 (n_12612, wc439, n_11947);
  not gc439 (wc439, n_12360);
  nand g28305 (n_12710, n_12405, n_12404);
  or g28306 (n_11864, n_11481, wc440);
  not gc440 (wc440, rst_n);
  nand g28307 (n_12112, rst_n, n_11469);
  or g28308 (n_12113, n_11469, wc441);
  not gc441 (wc441, rst_n);
  or g28309 (n_12601, n_11481, n_12599);
  nand g28311 (n_15340, n_12303, n_12302);
  nand g28312 (n_12772, n_12386, n_12385);
  nand g28313 (n_11812, n_12401, n_12400);
  nand g28314 (n_12766, n_12369, n_12368);
  nand g28316 (n_12703, n_12399, n_12398);
  or g28318 (n_12634, wc442, n_11950);
  not gc442 (wc442, n_11512);
  nand g28319 (n_11720, n_12389, n_12388);
  nand g28320 (n_11519, n_12371, n_12370);
  nand g28321 (n_12671, data_stack_pointer[1], n_11481);
  nand g28322 (n_12688, n_12373, n_12372);
  nand g28323 (n_12700, n_12393, n_12392);
  or g28324 (n_12172, n_11456, wc443);
  not gc443 (wc443, rst_n);
  or g28325 (n_12797, n_11456, n_12114);
  or g28326 (n_12153, \data_stack_mem[6] [7], n_11513);
  nand g28327 (n_12360, n_12538, n_11476);
  nand g28328 (n_12619, n_12384, n_12383);
  nand g28329 (n_12390, n_12120, n_12571);
  or g28330 (n_12386, \data_stack_mem[6] [1], n_11513);
  or g28331 (n_12395, \data_stack_mem[6] [4], n_11513);
  or g28332 (n_11950, sh_reg_in[8], wc444);
  not gc444 (wc444, n_12410);
  nand g28333 (n_12685, sh_reg_out_bit_counter[4], n_11455);
  nand g28334 (n_12622, n_12403, n_12402);
  or g28335 (n_12405, \data_stack_mem[6] [2], n_11513);
  nand g28336 (n_12388, n_12122, n_12568);
  or g28337 (n_12397, \data_stack_mem[6] [5], n_11513);
  nand g28338 (n_12400, n_12126, n_12574);
  nand g28340 (n_12370, n_11518, n_12562);
  or g28341 (n_12460, sh_reg_in[5], n_12459);
  or g28342 (n_12369, \data_stack_mem[6] [0], n_11513);
  or g28343 (n_12407, \data_stack_mem[6] [3], n_11513);
  nand g28344 (n_16359, n_12279, \data_stack_mem[0] [0]);
  or g28345 (n_16360, n_12279, \data_stack_mem[0] [0]);
  nand g28346 (n_11523, n_16359, n_16360);
  or g28347 (n_11575, n_12532, wc445);
  not gc445 (wc445, n_11508);
  nand g28349 (n_12380, n_12124, n_12565);
  nand g28350 (n_12507, sh_bit_cnt[3], n_11476);
  or g28351 (n_12377, \data_stack_mem[6] [6], n_11513);
  nand g28352 (n_12359, n_11455, n_12604);
  nand g28353 (n_11606, n_12531, n_15724);
  or g28356 (n_12459, sh_reg_in[7], n_12458);
  or g28357 (n_12571, wc446, n_11508);
  not gc446 (wc446, \data_stack_mem[0] [4]);
  or g28359 (n_12469, sh_reg_out_bit_counter[4], n_12468);
  or g28360 (n_12394, \data_stack_mem[5] [4], n_11515);
  nand g28361 (n_12532, n_12191, n_12531);
  or g28362 (n_12149, \data_stack_mem[5] [2], n_11515);
  or g28363 (n_12303, \data_stack_mem[5] [7], n_11515);
  or g28364 (n_12574, wc447, n_11508);
  not gc447 (wc447, \data_stack_mem[0] [7]);
  nand g28365 (n_12358, n_11454, n_12535);
  or g28366 (n_12562, wc448, n_11508);
  not gc448 (wc448, \data_stack_mem[0] [0]);
  nand g28367 (n_11513, n_11507, n_12330);
  or g28368 (n_12368, \data_stack_mem[5] [0], n_11515);
  nand g28369 (n_12604, sh_reg_out_bit_counter[3], n_11454);
  nand g28370 (n_12374, data_stack_pointer[3], n_12484);
  or g28371 (n_12565, wc449, n_11508);
  not gc449 (wc449, \data_stack_mem[0] [6]);
  or g28373 (n_12376, \data_stack_mem[5] [6], n_11515);
  nand g28374 (n_15724, \data_stack_mem[0] [1], n_12191);
  or g28375 (n_12385, \data_stack_mem[5] [1], n_11515);
  or g28376 (n_12568, wc450, n_11508);
  not gc450 (wc450, \data_stack_mem[0] [5]);
  or g28377 (n_12396, \data_stack_mem[5] [5], n_11515);
  or g28378 (n_12406, \data_stack_mem[5] [3], n_11515);
  nand g28379 (n_11504, data_stack_pointer[3], n_12496);
  nand g28380 (n_11947, n_12364, rst_n);
  or g28381 (n_11476, sh_bit_cnt[2], n_12480);
  nand g28382 (n_12332, n_11514, n_12472);
  or g28383 (n_11468, n_12419, wc451);
  not gc451 (wc451, rst_n);
  nand g28384 (n_12363, n_12480, n_12481);
  nand g28385 (n_11516, n_11507, n_12499);
  or g28386 (n_11517, wc452, n_11507);
  not gc452 (wc452, n_11512);
  or g28387 (n_12458, sh_reg_in[1], n_12457);
  or g28390 (n_12404, \data_stack_mem[3] [2], wc453);
  not gc453 (wc453, n_11507);
  or g28391 (n_12398, \data_stack_mem[3] [7], wc454);
  not gc454 (wc454, n_11507);
  or g28392 (n_12372, \data_stack_mem[3] [0], wc455);
  not gc455 (wc455, n_11507);
  or g28393 (n_12484, wc456, n_11503);
  not gc456 (wc456, \data_stack_mem[7] [0]);
  or g28394 (n_12378, \data_stack_mem[3] [6], wc457);
  not gc457 (wc457, n_11507);
  or g28395 (n_12392, \data_stack_mem[3] [5], wc458);
  not gc458 (wc458, n_11507);
  or g28396 (n_12496, data_stack_pointer[0], n_11503);
  nand g28397 (n_11496, n_11495, rst_n);
  or g28398 (n_12472, data_stack_pointer[1], wc459);
  not gc459 (wc459, n_12331);
  or g28399 (n_11882, data_stack_pointer[3], n_11881);
  or g28400 (n_12480, n_11475, enable_n);
  nand g28401 (n_12445, n_12442, n_12443);
  or g28403 (n_12468, sh_reg_out_bit_counter[3], n_12467);
  or g28404 (n_12531, wc460, n_11518);
  not gc460 (wc460, \data_stack_mem[1] [1]);
  or g28405 (n_12487, wc461, n_11503);
  not gc461 (wc461, data_stack_pointer[0]);
  nand g28406 (n_12361, n_11453, n_12475);
  or g28407 (n_12364, sh_bit_cnt[2], n_12448);
  nand g28408 (n_12419, n_12417, n_12418);
  or g28409 (n_12519, n_11862, wc462);
  not gc462 (wc462, rst_n);
  nand g28410 (n_12535, sh_reg_out_bit_counter[2], n_11453);
  nand g28411 (n_12538, sh_bit_cnt[2], n_11475);
  or g28412 (n_12559, n_12557, wc463);
  not gc463 (wc463, rst_n);
  nand g28413 (n_12261, \data_stack_mem[3] [0], n_11507);
  or g28414 (n_12499, data_stack_pointer[0], n_11514);
  or g28415 (n_11508, data_stack_pointer[1], n_11507);
  or g28416 (n_12599, n_11512, n_11968);
  or g28417 (n_12613, n_12611, wc464);
  not gc464 (wc464, rst_n);
  nand g28418 (n_12844, n_11538, rst_n);
  nand g28419 (n_12847, n_11546, rst_n);
  nand g28420 (n_12850, n_11532, rst_n);
  or g28421 (n_12882, data_stack_pointer[2], n_11485);
  nand g28422 (n_11515, n_11507, n_11514);
  or g28423 (n_13104, wc465, n_11485);
  not gc465 (wc465, data_stack_pointer[3]);
  or g28424 (n_11507, data_stack_pointer[2], data_stack_pointer[3]);
  nand g28425 (n_12120, \data_stack_mem[1] [4], \data_stack_mem[0] [4]);
  nand g28426 (n_12122, \data_stack_mem[1] [5], \data_stack_mem[0] [5]);
  nand g28427 (n_12124, \data_stack_mem[1] [6], \data_stack_mem[0] [6]);
  nand g28428 (n_12126, \data_stack_mem[1] [7], \data_stack_mem[0] [7]);
  or g28429 (n_12457, sh_reg_in[3], sh_reg_in[2]);
  or g28430 (n_11861, wc466, out_fifo_read_pointer[1]);
  not gc466 (wc466, out_fifo_read_pointer[0]);
  or g28431 (n_11862, out_fifo_read_pointer[0], wc467);
  not gc467 (wc467, out_fifo_read_pointer[1]);
  nand g28432 (n_11495, out_fifo_write_pointer[0],
       out_fifo_write_pointer[1]);
  or g28433 (n_11485, data_stack_pointer[0], wc468);
  not gc468 (wc468, rst_n);
  nand g28434 (n_11881, data_stack_pointer[0], rst_n);
  or g28435 (n_12444, wc469, out_fifo_write_pointer[0]);
  not gc469 (wc469, out_fifo_read_pointer[0]);
  or g28436 (n_12442, out_fifo_read_pointer[0], wc470);
  not gc470 (wc470, out_fifo_write_pointer[0]);
  or g28437 (n_12443, wc471, out_fifo_write_pointer[2]);
  not gc471 (wc471, out_fifo_read_pointer[2]);
  or g28438 (n_16361, wc472, out_fifo_write_pointer[1]);
  not gc472 (wc472, out_fifo_read_pointer[1]);
  or g28439 (n_16362, out_fifo_read_pointer[1], wc473);
  not gc473 (wc473, out_fifo_write_pointer[1]);
  nand g28440 (n_12441, n_16361, n_16362);
  nand g28441 (n_12114, rst_n, out_fifo_write_pointer[2]);
  or g28442 (n_12467, sh_reg_out_bit_counter[1],
       sh_reg_out_bit_counter[2]);
  nand g28443 (n_12781, data_stack_pointer[2], data_stack_pointer[3]);
  nand g28444 (n_12475, sh_reg_out_bit_counter[0],
       sh_reg_out_bit_counter[1]);
  or g28445 (n_12448, sh_bit_cnt[3], sh_bit_cnt[1]);
  or g28446 (n_12417, sh_bit_cnt[0], enable_n);
  nand g28447 (n_12418, sh_bit_cnt[0], enable_n);
  nand g28448 (n_12481, sh_bit_cnt[0], sh_bit_cnt[1]);
  nand g28449 (n_12557, sh_bit_cnt[1], enable_n);
  or g28450 (n_12592, data_stack_pointer[0], wc474);
  not gc474 (wc474, data_stack_pointer[1]);
  or g28451 (n_12590, wc475, data_stack_pointer[1]);
  not gc475 (wc475, data_stack_pointer[0]);
  or g28452 (n_12600, data_stack_pointer[2], wc476);
  not gc476 (wc476, data_stack_pointer[3]);
  nand g28453 (n_12611, sh_bit_cnt[2], enable_n);
  or g28454 (n_13099, data_stack_pointer[3], wc477);
  not gc477 (wc477, rst_n);
  or g28471 (n_11923, wc478, n_11922);
  not gc478 (wc478, n_12245);
  or g28472 (n_11924, wc479, n_11923);
  not gc479 (wc479, n_12186);
  or g28474 (n_12138, wc480, \data_stack_mem[3] [1]);
  not gc480 (wc480, n_11507);
  or g28475 (n_12148, wc481, \data_stack_mem[3] [3]);
  not gc481 (wc481, n_11507);
  or g28476 (n_12152, wc482, \data_stack_mem[3] [4]);
  not gc482 (wc482, n_11507);
  or g28477 (n_12231, n_11515, wc483);
  not gc483 (wc483, \data_stack_mem[5] [0]);
  or g28478 (n_12440, wc484, n_12445);
  not gc484 (wc484, n_12444);
  or g28479 (n_12410, n_12487, wc485);
  not gc485 (wc485, data_stack_pointer[3]);
  or g28480 (n_12197, n_11513, wc486);
  not gc486 (wc486, \data_stack_mem[6] [0]);
  or g28481 (n_11469, n_12469, wc487);
  not gc487 (wc487, sh_reg_out_bit_counter[0]);
  or g28482 (n_12558, wc488, n_11947);
  not gc488 (wc488, n_12363);
  or g28483 (n_11619, n_12622, wc489);
  not gc489 (wc489, \data_stack_mem[0] [2]);
  or g28484 (n_11585, n_12619, wc490);
  not gc490 (wc490, \data_stack_mem[0] [1]);
  or g28485 (n_12175, wc491, n_11950);
  not gc491 (wc491, rst_n);
  or g28487 (n_12583, n_11881, wc492);
  not gc492 (wc492, n_11481);
  or g28488 (n_12490, n_11501, wc493);
  not gc493 (wc493, sh_reg_in[0]);
  or g28489 (n_12718, n_11864, wc494);
  not gc494 (wc494, sh_reg_in[8]);
  or g28490 (n_12859, wc495, n_11457);
  not gc495 (wc495, n_12359);
  or g28491 (n_12856, wc496, n_11457);
  not gc496 (wc496, n_12358);
  or g28492 (n_12853, n_11457, n_12685);
  and g28493 (n_16342, wc497, sh_reg_out[21]);
  not gc497 (wc497, n_11457);
  and g28494 (n_16343, wc498, sh_reg_out[22]);
  not gc498 (wc498, n_11457);
  and g28495 (n_16344, wc499, sh_reg_out[23]);
  not gc499 (wc499, n_11457);
  and g28496 (n_16345, wc500, sh_reg_out[24]);
  not gc500 (wc500, n_11457);
  and g28497 (n_16346, wc501, sh_reg_out[8]);
  not gc501 (wc501, n_11457);
  and g28498 (n_16347, wc502, sh_reg_out[18]);
  not gc502 (wc502, n_11457);
  and g28499 (n_16348, wc503, sh_reg_out[25]);
  not gc503 (wc503, n_11457);
  and g28500 (n_16349, n_12361, wc504);
  not gc504 (wc504, n_11457);
  and g28501 (n_16350, wc505, sh_reg_out[26]);
  not gc505 (wc505, n_11457);
  and g28502 (n_16351, wc506, sh_reg_out[17]);
  not gc506 (wc506, n_11457);
  and g28503 (n_16352, wc507, sh_reg_out[16]);
  not gc507 (wc507, n_11457);
  and g28504 (n_16353, wc508, sh_reg_out[15]);
  not gc508 (wc508, n_11457);
  and g28505 (n_16354, wc509, sh_reg_out[14]);
  not gc509 (wc509, n_11457);
  or g28506 (n_11502, n_12493, wc510);
  not gc510 (wc510, sh_reg_in[4]);
  or g28507 (n_12712, n_12711, wc511);
  not gc511 (wc511, n_12147);
  or g28508 (n_12631, n_12630, wc512);
  not gc512 (wc512, n_12133);
  or g28509 (n_12786, wc513, n_11865);
  not gc513 (wc513, n_12332);
  or g28510 (n_11970, wc514, n_11482);
  not gc514 (wc514, n_12781);
  or g28511 (n_11621, n_12712, wc515);
  not gc515 (wc515, n_12149);
  or g28512 (n_11654, n_12631, wc516);
  not gc516 (wc516, \data_stack_mem[0] [3]);
  or g28513 (n_12871, n_11868, wc517);
  not gc517 (wc517, n_11968);
  or g28514 (n_12868, wc518, n_11868);
  not gc518 (wc518, n_11507);
  or g28515 (n_11908, n_12118, wc519);
  not gc519 (wc519, out_fifo_write_pointer[2]);
  or g28516 (n_11863, wc520, n_12520);
  not gc520 (wc520, n_12519);
  or g28517 (n_11563, n_12637, wc521);
  not gc521 (wc521, n_11509);
  or g28518 (n_11511, n_12640, wc522);
  not gc522 (wc522, n_11509);
  or g28519 (n_11981, wc523, n_11869);
  not gc523 (wc523, n_12871);
  or g28520 (n_11870, wc524, n_11869);
  not gc524 (wc524, n_12868);
  or g28521 (n_11486, n_12874, wc525);
  not gc525 (wc525, data_stack_pointer[3]);
  or g28522 (n_12841, wc526, n_12839);
  not gc526 (wc526, n_11507);
  or g28523 (n_11991, n_11981, wc527);
  not gc527 (wc527, n_11871);
  or g28524 (n_11982, n_11981, wc528);
  not gc528 (wc528, n_11866);
  or g28525 (n_11895, wc529, n_13105);
  not gc529 (wc529, n_11882);
  or g28526 (n_11913, n_11870, wc530);
  not gc530 (wc530, n_11866);
  or g28527 (n_12043, wc531, n_12883);
  not gc531 (wc531, n_11882);
  or g28528 (n_11872, n_11870, wc532);
  not gc532 (wc532, n_11871);
  or g28529 (n_13092, n_11577, wc533);
  not gc533 (wc533, n_12305);
  or g28530 (n_13093, wc534, n_12305);
  not gc534 (wc534, n_11577);
  or g28531 (n_13736, wc535, n_13732);
  not gc535 (wc535, n_13731);
  or g28532 (n_13688, wc536, n_13684);
  not gc536 (wc536, n_13683);
  or g28533 (n_14120, wc537, n_14116);
  not gc537 (wc537, n_14115);
  or g28534 (n_13976, wc538, n_13972);
  not gc538 (wc538, n_13971);
  or g28535 (n_13784, wc539, n_13780);
  not gc539 (wc539, n_13779);
  or g28536 (n_13640, wc540, n_13636);
  not gc540 (wc540, n_13635);
  or g28537 (n_14072, wc541, n_14068);
  not gc541 (wc541, n_14067);
  or g28538 (n_13496, wc542, n_13492);
  not gc542 (wc542, n_13491);
  or g28539 (n_13832, wc543, n_13828);
  not gc543 (wc543, n_13827);
  or g28540 (n_14264, wc544, n_14260);
  not gc544 (wc544, n_14259);
  or g28541 (n_13592, wc545, n_13588);
  not gc545 (wc545, n_13587);
  or g28542 (n_14168, wc546, n_14164);
  not gc546 (wc546, n_14163);
  or g28543 (n_13928, wc547, n_13924);
  not gc547 (wc547, n_13923);
  or g28544 (n_14024, wc548, n_14020);
  not gc548 (wc548, n_14019);
  or g28545 (n_13880, wc549, n_13876);
  not gc549 (wc549, n_13875);
  or g28546 (n_13544, wc550, n_13540);
  not gc550 (wc550, n_13539);
  or g28547 (n_14216, wc551, n_14212);
  not gc551 (wc551, n_14211);
  or g28548 (n_11603, wc552, n_14317);
  not gc552 (wc552, n_11507);
  or g28549 (n_14494, n_12148, wc553);
  not gc553 (wc553, n_11641);
  or g28550 (n_14493, wc554, n_14492);
  not gc554 (wc554, n_11507);
  or g28551 (n_11567, n_14476, wc555);
  not gc555 (wc555, data_stack_pointer[3]);
  or g28552 (n_12366, wc556, n_14470);
  not gc556 (wc556, n_14469);
  or g28553 (n_12287, wc557, n_14653);
  not gc557 (wc557, n_11507);
  or g28554 (n_14692, n_11505, wc558);
  not gc558 (wc558, n_11582);
  or g28555 (n_11598, n_14641, wc559);
  not gc559 (wc559, data_stack_pointer[3]);
  or g28556 (n_14539, n_11549, wc560);
  not gc560 (wc560, n_11530);
  or g28557 (n_14533, n_11541, wc561);
  not gc561 (wc561, n_11530);
  or g28558 (n_14527, n_11536, wc562);
  not gc562 (wc562, n_11530);
  or g28559 (n_14545, n_11553, wc563);
  not gc563 (wc563, n_11530);
  or g28560 (n_14551, n_11557, wc564);
  not gc564 (wc564, n_11530);
  or g28561 (n_14556, n_11561, wc565);
  not gc565 (wc565, n_11530);
  or g28562 (n_14569, n_11500, wc566);
  not gc566 (wc566, n_11530);
  or g28563 (n_14575, n_11544, wc567);
  not gc567 (wc567, n_11530);
  or g28564 (n_11705, wc568, n_14680);
  not gc568 (wc568, n_11507);
  or g28565 (n_14803, n_11769, wc569);
  not gc569 (wc569, n_12255);
  or g28566 (n_16290, wc570, \data_stack_mem[8] [2]);
  not gc570 (wc570, n_11615);
  or g28567 (n_16291, n_11615, wc571);
  not gc571 (wc571, \data_stack_mem[8] [2]);
  or g28568 (n_14797, n_11505, wc572);
  not gc572 (wc572, n_11615);
  or g28569 (n_11741, wc573, n_14779);
  not gc573 (wc573, n_11507);
  or g28570 (n_11634, n_14704, wc574);
  not gc574 (wc574, data_stack_pointer[3]);
  or g28571 (n_16280, wc575, \data_stack_mem[8] [3]);
  not gc575 (wc575, n_11631);
  or g28572 (n_16281, n_11631, wc576);
  not gc576 (wc576, \data_stack_mem[8] [3]);
  or g28573 (n_14920, n_11770, wc577);
  not gc577 (wc577, n_12181);
  or g28574 (n_11588, wc578, n_14731);
  not gc578 (wc578, n_14730);
  or g28575 (n_11822, n_11781, wc579);
  not gc579 (wc579, n_11784);
  or g28576 (n_14825, wc580, n_11651);
  not gc580 (wc580, n_11632);
  or g28577 (n_12258, n_11516, wc581);
  not gc581 (wc581, n_14992);
  or g28578 (n_15025, n_11771, wc582);
  not gc582 (wc582, n_12265);
  or g28579 (n_11666, n_14899, wc583);
  not gc583 (wc583, data_stack_pointer[3]);
  or g28580 (n_11622, wc584, n_14857);
  not gc584 (wc584, n_14856);
  or g28581 (n_11820, n_11780, wc585);
  not gc585 (wc585, n_11785);
  or g28582 (n_12168, n_11820, wc586);
  not gc586 (wc586, n_11823);
  or g28583 (n_16248, wc587, \data_stack_mem[8] [4]);
  not gc587 (wc587, n_11682);
  or g28584 (n_16249, n_11682, wc588);
  not gc588 (wc588, \data_stack_mem[8] [4]);
  or g28585 (n_15043, n_11505, wc589);
  not gc589 (wc589, n_11682);
  or g28586 (n_11656, wc590, n_14935);
  not gc590 (wc590, n_14934);
  or g28587 (n_12227, n_11515, wc591);
  not gc591 (wc591, n_15046);
  or g28588 (n_15055, n_11772, wc592);
  not gc592 (wc592, n_12264);
  or g28589 (n_11699, n_15013, wc593);
  not gc593 (wc593, data_stack_pointer[3]);
  or g28590 (n_11819, n_11779, wc594);
  not gc594 (wc594, n_11786);
  or g28591 (n_12233, n_11819, wc595);
  not gc595 (wc595, n_11824);
  or g28592 (n_15139, n_12153, wc596);
  not gc596 (wc596, n_11774);
  or g28593 (n_16232, wc597, \data_stack_mem[8] [5]);
  not gc597 (wc597, n_11716);
  or g28594 (n_16233, n_11716, wc598);
  not gc598 (wc598, \data_stack_mem[8] [5]);
  or g28595 (n_15145, n_11505, wc599);
  not gc599 (wc599, n_11716);
  or g28596 (n_15157, n_11773, wc600);
  not gc600 (wc600, n_12243);
  or g28597 (n_11735, n_15052, wc601);
  not gc601 (wc601, data_stack_pointer[3]);
  or g28598 (n_11689, wc602, n_15082);
  not gc602 (wc602, n_15081);
  or g28599 (n_11818, n_11778, wc603);
  not gc603 (wc603, n_11787);
  or g28600 (n_15240, n_11773, wc604);
  not gc604 (wc604, n_12291);
  or g28601 (n_15241, wc605, n_12291);
  not gc605 (wc605, n_11773);
  or g28602 (n_16218, wc606, \data_stack_mem[8] [6]);
  not gc606 (wc606, n_11732);
  or g28603 (n_16219, n_11732, wc607);
  not gc607 (wc607, \data_stack_mem[8] [6]);
  or g28604 (n_12245, n_11818, wc608);
  not gc608 (wc608, n_11825);
  or g28605 (n_15233, wc609, n_11752);
  not gc609 (wc609, n_11733);
  or g28606 (n_11777, n_12202, wc610);
  not gc610 (wc610, n_15247);
  or g28607 (n_16210, wc611, \data_stack_mem[8] [7]);
  not gc611 (wc611, n_11792);
  or g28608 (n_16211, n_11792, wc612);
  not gc612 (wc612, \data_stack_mem[8] [7]);
  or g28609 (n_12186, n_11817, wc613);
  not gc613 (wc613, n_11826);
  or g28610 (n_11723, wc614, n_15178);
  not gc614 (wc614, n_15177);
  or g28611 (n_15413, n_11789, wc615);
  not gc615 (wc615, n_11793);
  or g28612 (n_11757, wc616, n_15262);
  not gc616 (wc616, n_15261);
  or g28613 (n_16200, wc617, n_11588);
  not gc617 (wc617, n_11757);
  or g28614 (n_16201, n_11757, wc618);
  not gc618 (wc618, n_11588);
  or g28615 (n_15406, wc619, n_11828);
  not gc619 (wc619, n_11924);
  or g28616 (n_11927, n_15406, wc620);
  not gc620 (wc620, n_11827);
  or g28617 (n_11815, wc621, n_15346);
  not gc621 (wc621, n_15345);
  or g28618 (n_15433, n_11549, wc622);
  not gc622 (wc622, n_11794);
  or g28619 (n_15427, n_11541, wc623);
  not gc623 (wc623, n_11794);
  or g28620 (n_15439, n_11553, wc624);
  not gc624 (wc624, n_11794);
  or g28621 (n_15421, n_11536, wc625);
  not gc625 (wc625, n_11794);
  or g28622 (n_15445, n_11557, wc626);
  not gc626 (wc626, n_11794);
  or g28623 (n_15511, n_11544, wc627);
  not gc627 (wc627, n_11794);
  or g28624 (n_15450, n_11561, wc628);
  not gc628 (wc628, n_11794);
  or g28625 (n_15505, n_11500, wc629);
  not gc629 (wc629, n_11794);
  or g28626 (n_12012, n_11830, wc630);
  not gc630 (wc630, n_11927);
  or g28627 (n_16190, wc631, n_11530);
  not gc631 (wc631, n_11815);
  or g28628 (n_16191, n_11815, wc632);
  not gc632 (wc632, n_11530);
  or g28629 (n_15526, n_11536, wc633);
  not gc633 (wc633, n_11830);
  or g28630 (n_15532, n_11541, wc634);
  not gc634 (wc634, n_11830);
  or g28631 (n_15538, n_11549, wc635);
  not gc635 (wc635, n_11830);
  or g28632 (n_15544, n_11553, wc636);
  not gc636 (wc636, n_11830);
  or g28633 (n_15550, n_11557, wc637);
  not gc637 (wc637, n_11830);
  or g28634 (n_15555, n_11561, wc638);
  not gc638 (wc638, n_11830);
  or g28635 (n_16182, wc639, n_11794);
  not gc639 (wc639, n_12012);
  or g28636 (n_16183, n_12012, wc640);
  not gc640 (wc640, n_11794);
  or g28637 (n_15631, n_11536, wc641);
  not gc641 (wc641, n_11925);
  or g28638 (n_15655, n_11557, wc642);
  not gc642 (wc642, n_11925);
  or g28639 (n_15649, n_11553, wc643);
  not gc643 (wc643, n_11925);
  or g28640 (n_15643, n_11549, wc644);
  not gc644 (wc644, n_11925);
  or g28641 (n_15673, n_11544, wc645);
  not gc645 (wc645, n_11925);
  or g28642 (n_15637, n_11541, wc646);
  not gc646 (wc646, n_11925);
  or g28643 (n_15667, n_11500, wc647);
  not gc647 (wc647, n_11925);
  or g28644 (n_15660, n_11561, wc648);
  not gc648 (wc648, n_11925);
  or g28645 (n_15703, n_11553, wc649);
  not gc649 (wc649, n_12014);
  or g28646 (n_15697, n_11549, wc650);
  not gc650 (wc650, n_12014);
  or g28647 (n_15714, n_11561, wc651);
  not gc651 (wc651, n_12014);
  or g28648 (n_15709, n_11557, wc652);
  not gc652 (wc652, n_12014);
  or g28649 (n_15685, n_11536, wc653);
  not gc653 (wc653, n_12014);
  or g28650 (n_15691, n_11541, wc654);
  not gc654 (wc654, n_12014);
  or g28651 (n_15586, n_11549, wc655);
  not gc655 (wc655, n_11852);
  or g28652 (n_15598, n_11557, wc656);
  not gc656 (wc656, n_11852);
  or g28653 (n_15574, n_11536, wc657);
  not gc657 (wc657, n_11852);
  or g28654 (n_15592, n_11553, wc658);
  not gc658 (wc658, n_11852);
  or g28655 (n_15580, n_11541, wc659);
  not gc659 (wc659, n_11852);
  or g28656 (n_15603, n_11561, wc660);
  not gc660 (wc660, n_11852);
  CDN_flop \out_fifo_read_pointer_reg[0] (.clk (clk), .d (n_11470),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[0]));
  CDN_flop \out_fifo_read_pointer_reg[1] (.clk (clk), .d (n_11863),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[1]));
  CDN_flop \out_fifo_read_pointer_reg[2] (.clk (clk), .d (n_12024),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[2]));
  CDN_flop \out_fifo_reg[0][0][0] (.clk (clk), .d (n_11854), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [0]));
  CDN_flop \out_fifo_reg[0][0][1] (.clk (clk), .d (n_11537), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [1]));
  CDN_flop \out_fifo_reg[0][0][2] (.clk (clk), .d (n_11590), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [2]));
  CDN_flop \out_fifo_reg[0][0][3] (.clk (clk), .d (n_11624), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [3]));
  CDN_flop \out_fifo_reg[0][0][4] (.clk (clk), .d (n_11658), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [4]));
  CDN_flop \out_fifo_reg[0][0][5] (.clk (clk), .d (n_11691), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [5]));
  CDN_flop \out_fifo_reg[0][0][6] (.clk (clk), .d (n_11725), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [6]));
  CDN_flop \out_fifo_reg[0][0][7] (.clk (clk), .d (n_11796), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [7]));
  CDN_flop \out_fifo_reg[0][0][8] (.clk (clk), .d (n_11832), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [8]));
  CDN_flop \out_fifo_reg[0][1][0] (.clk (clk), .d (n_12016), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [0]));
  CDN_flop \out_fifo_reg[0][1][1] (.clk (clk), .d (n_11797), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [1]));
  CDN_flop \out_fifo_reg[0][1][2] (.clk (clk), .d (n_11833), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [2]));
  CDN_flop \out_fifo_reg[0][1][3] (.clk (clk), .d (n_11929), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [3]));
  CDN_flop \out_fifo_reg[0][1][4] (.clk (clk), .d (n_11928), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [4]));
  CDN_flop \out_fifo_reg[0][2][0] (.clk (clk), .d (n_12036), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [0]));
  CDN_flop \out_fifo_reg[0][2][1] (.clk (clk), .d (n_12031), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [1]));
  CDN_flop \out_fifo_reg[0][2][8] (.clk (clk), .d (n_11959), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [8]));
  CDN_flop \out_fifo_reg[0][2][9] (.clk (clk), .d (1'b1), .sena
       (n_11945), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (\out_fifo[0][2] [9]));
  CDN_flop \out_fifo_reg[1][0][0] (.clk (clk), .d (n_11857), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [0]));
  CDN_flop \out_fifo_reg[1][0][1] (.clk (clk), .d (n_11550), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [1]));
  CDN_flop \out_fifo_reg[1][0][2] (.clk (clk), .d (n_11593), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [2]));
  CDN_flop \out_fifo_reg[1][0][3] (.clk (clk), .d (n_11627), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [3]));
  CDN_flop \out_fifo_reg[1][0][4] (.clk (clk), .d (n_11661), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [4]));
  CDN_flop \out_fifo_reg[1][0][5] (.clk (clk), .d (n_11694), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [5]));
  CDN_flop \out_fifo_reg[1][0][6] (.clk (clk), .d (n_11728), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [6]));
  CDN_flop \out_fifo_reg[1][0][7] (.clk (clk), .d (n_11802), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [7]));
  CDN_flop \out_fifo_reg[1][0][8] (.clk (clk), .d (n_11838), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [8]));
  CDN_flop \out_fifo_reg[1][1][0] (.clk (clk), .d (n_12019), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [0]));
  CDN_flop \out_fifo_reg[1][1][1] (.clk (clk), .d (n_11803), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [1]));
  CDN_flop \out_fifo_reg[1][1][2] (.clk (clk), .d (n_11839), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [2]));
  CDN_flop \out_fifo_reg[1][1][3] (.clk (clk), .d (n_11934), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [3]));
  CDN_flop \out_fifo_reg[1][1][4] (.clk (clk), .d (n_11933), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [4]));
  CDN_flop \out_fifo_reg[1][2][0] (.clk (clk), .d (n_12039), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [0]));
  CDN_flop \out_fifo_reg[1][2][1] (.clk (clk), .d (n_12030), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [1]));
  CDN_flop \out_fifo_reg[1][2][8] (.clk (clk), .d (n_11961), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [8]));
  CDN_flop \out_fifo_reg[1][2][9] (.clk (clk), .d (1'b1), .sena
       (n_11942), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (\out_fifo[1][2] [9]));
  CDN_flop \out_fifo_reg[2][0][0] (.clk (clk), .d (n_11858), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [0]));
  CDN_flop \out_fifo_reg[2][0][1] (.clk (clk), .d (n_11554), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [1]));
  CDN_flop \out_fifo_reg[2][0][2] (.clk (clk), .d (n_11594), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [2]));
  CDN_flop \out_fifo_reg[2][0][3] (.clk (clk), .d (n_11628), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [3]));
  CDN_flop \out_fifo_reg[2][0][4] (.clk (clk), .d (n_11662), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [4]));
  CDN_flop \out_fifo_reg[2][0][5] (.clk (clk), .d (n_11695), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [5]));
  CDN_flop \out_fifo_reg[2][0][6] (.clk (clk), .d (n_11729), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [6]));
  CDN_flop \out_fifo_reg[2][0][7] (.clk (clk), .d (n_11804), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [7]));
  CDN_flop \out_fifo_reg[2][0][8] (.clk (clk), .d (n_11840), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [8]));
  CDN_flop \out_fifo_reg[2][1][0] (.clk (clk), .d (n_12020), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [0]));
  CDN_flop \out_fifo_reg[2][1][1] (.clk (clk), .d (n_11805), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [1]));
  CDN_flop \out_fifo_reg[2][1][2] (.clk (clk), .d (n_11841), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [2]));
  CDN_flop \out_fifo_reg[2][1][3] (.clk (clk), .d (n_11936), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [3]));
  CDN_flop \out_fifo_reg[2][1][4] (.clk (clk), .d (n_11935), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [4]));
  CDN_flop \out_fifo_reg[2][2][0] (.clk (clk), .d (n_12040), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [0]));
  CDN_flop \out_fifo_reg[2][2][1] (.clk (clk), .d (n_12032), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [1]));
  CDN_flop \out_fifo_reg[2][2][8] (.clk (clk), .d (n_11962), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [8]));
  CDN_flop \out_fifo_reg[2][2][9] (.clk (clk), .d (1'b1), .sena
       (n_11943), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (\out_fifo[2][2] [9]));
  CDN_flop \out_fifo_reg[3][0][0] (.clk (clk), .d (n_11856), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [0]));
  CDN_flop \out_fifo_reg[3][0][1] (.clk (clk), .d (n_11545), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [1]));
  CDN_flop \out_fifo_reg[3][0][2] (.clk (clk), .d (n_11592), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [2]));
  CDN_flop \out_fifo_reg[3][0][3] (.clk (clk), .d (n_11626), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [3]));
  CDN_flop \out_fifo_reg[3][0][4] (.clk (clk), .d (n_11660), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [4]));
  CDN_flop \out_fifo_reg[3][0][5] (.clk (clk), .d (n_11693), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [5]));
  CDN_flop \out_fifo_reg[3][0][6] (.clk (clk), .d (n_11727), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [6]));
  CDN_flop \out_fifo_reg[3][0][7] (.clk (clk), .d (n_11800), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [7]));
  CDN_flop \out_fifo_reg[3][0][8] (.clk (clk), .d (n_11836), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [8]));
  CDN_flop \out_fifo_reg[3][1][0] (.clk (clk), .d (n_12018), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [0]));
  CDN_flop \out_fifo_reg[3][1][1] (.clk (clk), .d (n_11801), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [1]));
  CDN_flop \out_fifo_reg[3][1][2] (.clk (clk), .d (n_11837), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [2]));
  CDN_flop \out_fifo_reg[3][1][3] (.clk (clk), .d (n_11932), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [3]));
  CDN_flop \out_fifo_reg[3][1][4] (.clk (clk), .d (n_12011), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [4]));
  CDN_flop \out_fifo_reg[3][2][0] (.clk (clk), .d (n_12038), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [0]));
  CDN_flop \out_fifo_reg[3][2][1] (.clk (clk), .d (n_12033), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [1]));
  CDN_flop \out_fifo_reg[3][2][8] (.clk (clk), .d (n_11956), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [8]));
  CDN_flop \out_fifo_reg[3][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16337), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (\out_fifo[3][2] [9]));
  CDN_flop \out_fifo_reg[4][0][0] (.clk (clk), .d (n_11859), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [0]));
  CDN_flop \out_fifo_reg[4][0][1] (.clk (clk), .d (n_11558), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [1]));
  CDN_flop \out_fifo_reg[4][0][2] (.clk (clk), .d (n_11595), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [2]));
  CDN_flop \out_fifo_reg[4][0][3] (.clk (clk), .d (n_11629), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [3]));
  CDN_flop \out_fifo_reg[4][0][4] (.clk (clk), .d (n_11663), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [4]));
  CDN_flop \out_fifo_reg[4][0][5] (.clk (clk), .d (n_11696), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [5]));
  CDN_flop \out_fifo_reg[4][0][6] (.clk (clk), .d (n_11730), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [6]));
  CDN_flop \out_fifo_reg[4][0][7] (.clk (clk), .d (n_11806), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [7]));
  CDN_flop \out_fifo_reg[4][0][8] (.clk (clk), .d (n_11842), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [8]));
  CDN_flop \out_fifo_reg[4][1][0] (.clk (clk), .d (n_12021), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [0]));
  CDN_flop \out_fifo_reg[4][1][1] (.clk (clk), .d (n_11807), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [1]));
  CDN_flop \out_fifo_reg[4][1][2] (.clk (clk), .d (n_11843), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [2]));
  CDN_flop \out_fifo_reg[4][1][3] (.clk (clk), .d (n_11938), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [3]));
  CDN_flop \out_fifo_reg[4][1][4] (.clk (clk), .d (n_11937), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [4]));
  CDN_flop \out_fifo_reg[4][2][0] (.clk (clk), .d (n_12041), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [0]));
  CDN_flop \out_fifo_reg[4][2][1] (.clk (clk), .d (n_11911), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [1]));
  CDN_flop \out_fifo_reg[4][2][8] (.clk (clk), .d (n_11963), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [8]));
  CDN_flop \out_fifo_reg[4][2][9] (.clk (clk), .d (1'b1), .sena
       (n_11941), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (\out_fifo[4][2] [9]));
  CDN_flop \out_fifo_reg[5][0][0] (.clk (clk), .d (n_11860), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [0]));
  CDN_flop \out_fifo_reg[5][0][1] (.clk (clk), .d (n_11562), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [1]));
  CDN_flop \out_fifo_reg[5][0][2] (.clk (clk), .d (n_11596), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [2]));
  CDN_flop \out_fifo_reg[5][0][3] (.clk (clk), .d (n_11630), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [3]));
  CDN_flop \out_fifo_reg[5][0][4] (.clk (clk), .d (n_11664), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [4]));
  CDN_flop \out_fifo_reg[5][0][5] (.clk (clk), .d (n_11697), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [5]));
  CDN_flop \out_fifo_reg[5][0][6] (.clk (clk), .d (n_11731), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [6]));
  CDN_flop \out_fifo_reg[5][0][7] (.clk (clk), .d (n_11808), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [7]));
  CDN_flop \out_fifo_reg[5][0][8] (.clk (clk), .d (n_11844), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [8]));
  CDN_flop \out_fifo_reg[5][1][0] (.clk (clk), .d (n_12022), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [0]));
  CDN_flop \out_fifo_reg[5][1][1] (.clk (clk), .d (n_11809), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [1]));
  CDN_flop \out_fifo_reg[5][1][2] (.clk (clk), .d (n_11845), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [2]));
  CDN_flop \out_fifo_reg[5][1][3] (.clk (clk), .d (n_11940), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [3]));
  CDN_flop \out_fifo_reg[5][1][4] (.clk (clk), .d (n_11939), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [4]));
  CDN_flop \out_fifo_reg[5][2][0] (.clk (clk), .d (n_12042), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [0]));
  CDN_flop \out_fifo_reg[5][2][1] (.clk (clk), .d (n_11909), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [1]));
  CDN_flop \out_fifo_reg[5][2][8] (.clk (clk), .d (n_11964), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [8]));
  CDN_flop \out_fifo_reg[5][2][9] (.clk (clk), .d (1'b1), .sena
       (n_11944), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (\out_fifo[5][2] [9]));
  CDN_flop \out_fifo_reg[6][0][0] (.clk (clk), .d (n_11855), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [0]));
  CDN_flop \out_fifo_reg[6][0][1] (.clk (clk), .d (n_11542), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [1]));
  CDN_flop \out_fifo_reg[6][0][2] (.clk (clk), .d (n_11591), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [2]));
  CDN_flop \out_fifo_reg[6][0][3] (.clk (clk), .d (n_11625), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [3]));
  CDN_flop \out_fifo_reg[6][0][4] (.clk (clk), .d (n_11659), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [4]));
  CDN_flop \out_fifo_reg[6][0][5] (.clk (clk), .d (n_11692), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [5]));
  CDN_flop \out_fifo_reg[6][0][6] (.clk (clk), .d (n_11726), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [6]));
  CDN_flop \out_fifo_reg[6][0][7] (.clk (clk), .d (n_11798), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [7]));
  CDN_flop \out_fifo_reg[6][0][8] (.clk (clk), .d (n_11834), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [8]));
  CDN_flop \out_fifo_reg[6][1][0] (.clk (clk), .d (n_12017), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [0]));
  CDN_flop \out_fifo_reg[6][1][1] (.clk (clk), .d (n_11799), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [1]));
  CDN_flop \out_fifo_reg[6][1][2] (.clk (clk), .d (n_11835), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [2]));
  CDN_flop \out_fifo_reg[6][1][3] (.clk (clk), .d (n_11931), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [3]));
  CDN_flop \out_fifo_reg[6][1][4] (.clk (clk), .d (n_11930), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [4]));
  CDN_flop \out_fifo_reg[6][2][0] (.clk (clk), .d (n_12037), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [0]));
  CDN_flop \out_fifo_reg[6][2][1] (.clk (clk), .d (n_11910), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [1]));
  CDN_flop \out_fifo_reg[6][2][8] (.clk (clk), .d (n_11960), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [8]));
  CDN_flop \out_fifo_reg[6][2][9] (.clk (clk), .d (1'b1), .sena
       (n_11946), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (\out_fifo[6][2] [9]));
  CDN_flop \out_fifo_reg[7][0][0] (.clk (clk), .d (n_11853), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [0]));
  CDN_flop \out_fifo_reg[7][0][1] (.clk (clk), .d (n_11531), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [1]));
  CDN_flop \out_fifo_reg[7][0][2] (.clk (clk), .d (n_11589), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [2]));
  CDN_flop \out_fifo_reg[7][0][3] (.clk (clk), .d (n_11623), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [3]));
  CDN_flop \out_fifo_reg[7][0][4] (.clk (clk), .d (n_11657), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [4]));
  CDN_flop \out_fifo_reg[7][0][5] (.clk (clk), .d (n_11690), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [5]));
  CDN_flop \out_fifo_reg[7][0][6] (.clk (clk), .d (n_11724), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [6]));
  CDN_flop \out_fifo_reg[7][0][7] (.clk (clk), .d (n_11758), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [7]));
  CDN_flop \out_fifo_reg[7][0][8] (.clk (clk), .d (n_11816), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [8]));
  CDN_flop \out_fifo_reg[7][1][0] (.clk (clk), .d (n_12015), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [0]));
  CDN_flop \out_fifo_reg[7][1][1] (.clk (clk), .d (n_11795), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [1]));
  CDN_flop \out_fifo_reg[7][1][2] (.clk (clk), .d (n_11831), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [2]));
  CDN_flop \out_fifo_reg[7][1][3] (.clk (clk), .d (n_11926), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [3]));
  CDN_flop \out_fifo_reg[7][1][4] (.clk (clk), .d (n_12010), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [4]));
  CDN_flop \out_fifo_reg[7][2][0] (.clk (clk), .d (n_12035), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [0]));
  CDN_flop \out_fifo_reg[7][2][1] (.clk (clk), .d (n_11958), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [1]));
  CDN_flop \out_fifo_reg[7][2][8] (.clk (clk), .d (n_11955), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [8]));
  CDN_flop \out_fifo_reg[7][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16336), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (\out_fifo[7][2] [9]));
  CDN_flop \out_fifo_write_pointer_reg[0] (.clk (clk), .d (n_11953),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[0]));
  CDN_flop \out_fifo_write_pointer_reg[1] (.clk (clk), .d (n_11954),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[1]));
  CDN_flop \out_fifo_write_pointer_reg[2] (.clk (clk), .d (n_12023),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[2]));
  CDN_flop \sh_bit_cnt_reg[0] (.clk (clk), .d (n_11468), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[0]));
  CDN_flop \sh_bit_cnt_reg[1] (.clk (clk), .d (n_11949), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[1]));
  CDN_flop \sh_bit_cnt_reg[2] (.clk (clk), .d (n_11948), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[2]));
  CDN_flop \sh_bit_cnt_reg[3] (.clk (clk), .d (n_11477), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[3]));
  CDN_flop \sh_reg_in_reg[0] (.clk (clk), .d (din), .sena (n_11463),
       .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd (1'b0), .q
       (sh_reg_in[0]));
  CDN_flop \sh_reg_in_reg[1] (.clk (clk), .d (sh_reg_in[0]), .sena
       (n_11463), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (sh_reg_in[1]));
  CDN_flop \sh_reg_in_reg[2] (.clk (clk), .d (sh_reg_in[1]), .sena
       (n_11463), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (sh_reg_in[2]));
  CDN_flop \sh_reg_in_reg[3] (.clk (clk), .d (sh_reg_in[2]), .sena
       (n_11463), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (sh_reg_in[3]));
  CDN_flop \sh_reg_in_reg[4] (.clk (clk), .d (sh_reg_in[3]), .sena
       (n_11463), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (sh_reg_in[4]));
  CDN_flop \sh_reg_in_reg[5] (.clk (clk), .d (sh_reg_in[4]), .sena
       (n_11463), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (sh_reg_in[5]));
  CDN_flop \sh_reg_in_reg[6] (.clk (clk), .d (sh_reg_in[5]), .sena
       (n_11463), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (sh_reg_in[6]));
  CDN_flop \sh_reg_in_reg[7] (.clk (clk), .d (sh_reg_in[6]), .sena
       (n_11463), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (sh_reg_in[7]));
  CDN_flop \sh_reg_in_reg[8] (.clk (clk), .d (sh_reg_in[7]), .sena
       (n_11463), .aclr (1'b0), .apre (1'b0), .srl (n_11462), .srd
       (1'b0), .q (sh_reg_in[8]));
  CDN_flop \sh_reg_out_bit_counter_reg[0] (.clk (clk), .d (n_11480),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[0]));
  CDN_flop \sh_reg_out_bit_counter_reg[1] (.clk (clk), .d (n_16349),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[1]));
  CDN_flop \sh_reg_out_bit_counter_reg[2] (.clk (clk), .d (n_11967),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[2]));
  CDN_flop \sh_reg_out_bit_counter_reg[3] (.clk (clk), .d (n_11966),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[3]));
  CDN_flop \sh_reg_out_bit_counter_reg[4] (.clk (clk), .d (n_11965),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[4]));
  CDN_flop \sh_reg_out_reg[0] (.clk (clk), .d (n_12009), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[0]));
  CDN_flop \sh_reg_out_reg[1] (.clk (clk), .d (n_12065), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[1]));
  CDN_flop \sh_reg_out_reg[2] (.clk (clk), .d (n_12064), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[2]));
  CDN_flop \sh_reg_out_reg[3] (.clk (clk), .d (n_12063), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[3]));
  CDN_flop \sh_reg_out_reg[4] (.clk (clk), .d (n_12062), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[4]));
  CDN_flop \sh_reg_out_reg[5] (.clk (clk), .d (n_12060), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[5]));
  CDN_flop \sh_reg_out_reg[6] (.clk (clk), .d (n_12059), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[6]));
  CDN_flop \sh_reg_out_reg[7] (.clk (clk), .d (n_12061), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[7]));
  CDN_flop \sh_reg_out_reg[8] (.clk (clk), .d (n_12057), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[8]));
  CDN_flop \sh_reg_out_reg[9] (.clk (clk), .d (n_16346), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[9]));
  CDN_flop \sh_reg_out_reg[10] (.clk (clk), .d (n_12066), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[10]));
  CDN_flop \sh_reg_out_reg[11] (.clk (clk), .d (n_12056), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[11]));
  CDN_flop \sh_reg_out_reg[12] (.clk (clk), .d (n_12054), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[12]));
  CDN_flop \sh_reg_out_reg[13] (.clk (clk), .d (n_12053), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[13]));
  CDN_flop \sh_reg_out_reg[14] (.clk (clk), .d (n_12068), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[14]));
  CDN_flop \sh_reg_out_reg[15] (.clk (clk), .d (n_16354), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[15]));
  CDN_flop \sh_reg_out_reg[16] (.clk (clk), .d (n_16353), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[16]));
  CDN_flop \sh_reg_out_reg[17] (.clk (clk), .d (n_16352), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[17]));
  CDN_flop \sh_reg_out_reg[18] (.clk (clk), .d (n_16351), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[18]));
  CDN_flop \sh_reg_out_reg[19] (.clk (clk), .d (n_16347), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[19]));
  CDN_flop \sh_reg_out_reg[20] (.clk (clk), .d (n_12067), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[20]));
  CDN_flop \sh_reg_out_reg[21] (.clk (clk), .d (n_12069), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[21]));
  CDN_flop \sh_reg_out_reg[22] (.clk (clk), .d (n_16342), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[22]));
  CDN_flop \sh_reg_out_reg[23] (.clk (clk), .d (n_16343), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[23]));
  CDN_flop \sh_reg_out_reg[24] (.clk (clk), .d (n_16344), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[24]));
  CDN_flop \sh_reg_out_reg[25] (.clk (clk), .d (n_16345), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[25]));
  CDN_flop \sh_reg_out_reg[26] (.clk (clk), .d (n_16348), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[26]));
  CDN_flop \sh_reg_out_reg[27] (.clk (clk), .d (n_16350), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[27]));
  CDN_flop \sh_reg_out_reg[28] (.clk (clk), .d (n_12058), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[28]));
  CDN_flop \sh_reg_out_reg[29] (.clk (clk), .d (n_12055), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (dout));
endmodule

`ifdef RC_CDN_GENERIC_GATE
`else
module CDN_flop(clk, d, sena, aclr, apre, srl, srd, q);
  input clk, d, sena, aclr, apre, srl, srd;
  output q;
  wire clk, d, sena, aclr, apre, srl, srd;
  wire q;
  reg  qi;
  assign #1 q = qi;
  always 
    @(posedge clk or posedge apre or posedge aclr) 
      if (aclr) 
        qi <= 0;
      else if (apre) 
          qi <= 1;
        else if (srl) 
            qi <= srd;
          else begin
            if (sena) 
              qi <= d;
          end
  initial 
    qi <= 1'b0;
endmodule
`endif
