/******************************************************************************
 * (C) Copyright 2022 AGH UST All Rights Reserved
 ******************************************************************************
 * MODULE NAME: vdic_dut_2022
 * VERSION:     1.4
 * DATE:        01-12-2022
 *
 * ABSTRACT:   DUT module for VDIC 2022 labs.
 *              The DUT is RPN calculator type. The arguments are sent first,
 *              than the operator/command.
 *******************************************************************************
 * HISTORY:
 * 20-10-2022 v1.0 Initial version
 * 03-11-2022 v1.1 Added remaining commands
 * 10-11-2022 v1.2 Modifications:
 *            - corrected bug: zero returned for invalid command
 *            - corrected spec: CMD_AND description
 * 24-11-2022 v1.3 Modifications:
 *            - corrected operation for 10 args
 *            - implemented data parity checking
 * 01-12-2022 v1.4 Modifications:
 *            - implemented command parity checking
 * 
 *******************************************************************************
 * INPUTS
 *    clk      - posedge active clock, always running
 *    rst_n    - synchronous reset active low
 *    din      - serial data input
 *    enable_n - chip enable, active low;

 * OUTPUTS
 *    dout       - serial data output
 *    dout_valid - valid flag for serial data output, active high
 *
 *******************************************************************************

 The clock is always active.
 The DUT operates on the posedge of the clock.
 The DUT receives the data when enable_n is active.
 IMPORTANT: din and dout can operate in parallel - DUT has some internal buffering
 implemented.

 --------------------------------------------------------------------------------
 --- Input data
 --------------------------------------------------------------------------------

 The input data is send serially in WORDs.

 The WORD is always 10 bit long. MSB is sent first.
 The WORD sent to the DUT is either DATA type or CONTROL type.

 DATA = 0bbbbbbbbp
 where:
 - b = 0 or 1, PAYLOAD bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 CONTROL = 1bbbbbbbbp
 where:
 - b = 0 or 1, COMMAND bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 The COMMAND can be:
 00000000 - CMD_NOP, do nothing, remove the data (reset data stack)
 00000001 - CMD_AND, logic AND of the arguments
 00000010 - CMD_OR, logic OR of the arguments
 00000011 - CMD_XOR, logic XOR of the arguments
 00010000 - CMD_ADD, add the arguments
 00100000 - CMD_SUB, subtract other arguments from the first one

 --------------------------------------------------------------------------------
 --- Output data
 --------------------------------------------------------------------------------

 The DUT responds to each CONTROL word, sending 3 WORDS:
 STATUS, DATA, DATA

 STATUS = 1bbbbbbbbp
 where bbbbbbbb is one of:

 00000000 - S_NO_ERROR - data correctly processed
 00000001 - S_MISSING_DATA - missing input data
 00000010 - S_DATA_STACK_OVERFLOW - maximum number of arguments exceeded
 00000100 - S_OUTPUT_FIFO_OVERFLOW - result dropped not possible to process
 00100000 - S_DATA_PARITY_ERROR - input data or command parity error
 01000000 - S_COMMAND_PARITY_ERROR - input data or command parity error
 10000000 - S_INVALID_COMMAND - unknown command detected

 DATA is defined as in the input.
 PAYLOAD of the DATA is 00000000 if the data was NOT processed correctly.

 *******************************************************************************
 * IMPLEMENTATION STATUS
 *******************************************************************************
 *  <Feature>                        <Is implemented>
 *    command CMD_NOP                   YES
 *    command CMD_AND                   YES
 *    command CMD_OR                    YES
 *    command CMD_XOR                   YES
 *    command CMD_ADD                   YES
 *    command CMD_SUB                   YES
 *    status S_NO_ERROR                 YES
 *    status S_MISSING_DATA              NO
 *    status S_DATA_STACK_OVERFLOW       NO
 *    status S_OUTPUT_FIFO_OVERFLOW      NO
 *    status S_DATA_PARITY_ERROR        YES
 *    status S_COMMAND_PARITY_ERROR     YES
 *    status S_INVALID_COMMAND          YES
 *******************************************************************************
 */
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
jONIetVf9Mdyg/iVn4m1+IYRHWWBErqo9Sf3/82cc8+I65YN6316vwJsLMph52rq
2o2uRDqgb9J97wP2YTJnCDEYgOtPLheXlMKPwRhSsKVkiCyYXfQA/34naZ5AafYB
MURChIrP0c5h+DTXRzzZbJp9KVBr77KGmeEBpH5jq2Fnj3tOGcfOG9gxGH8XohmA
EOytr08jfMQZr+F1cLeq2XqmvVKOJA9aWkU+KUBaKd7Yi8N2yeq32bHLPq1sOJ8A
rzt36UAICH2rA7jeKb0VNmlLE4i88qQ265dbPCMAE6cd3hXiXmA/TSKuwybomkHa
72uJAyNjcOfBxE8BchKmeA==
//pragma protect end_key_block
//pragma protect digest_block
7g7oJoE2R1VUIBQ7/7vOpPox93U=
//pragma protect end_digest_block
//pragma protect data_block
rluRA5rd3YH2lbZYLfBdVOYPGZdkBY23QS1o7vO9z3pEca/r1xdfmQDE2WXxEMjZ
quqA3DT+p7YFrKy9rJyv+rE4nmxUZmFl4tFEEUd+B4E5VK2mds2jYO5ECWChzKn1
FFlYIT+jdkrffSJOFFcXAOxGI76q586pufmf+Dop24BgOq50n4AmDC558HwLiTvz
Y/4uGZLmu+C5qy9PWdrfKDqM4XsButv7fAbjJzr2JfZvAvGU2aM1jTiAEBx9t+ad
jqV78/RlHeDzWAJrdskTm7MryL8INEAQ/TUHeXYwjtoQlGXcDjeE3q9f39DNRxVd
dJUjLNb2LPETgE073AY3T8RN81PIS1UFe4w9yiD2/1mSy3TLtptUwnarKT/CQiyl
CmxLEgdnbDk1nw+cGzqQZ5+Q3hdKStMxaHYxyNyhF4e40IZv7Xd5LfHaIEOjd5OC
S30SqivaAm22E+cr0PdjcuNnimBYY+s6+jE5/XAUQ1mfs0LdM8JMiJEp6dgWkohD
tTxjsaW1liwuf/ifn4Yh0IQTBYHyTD24QYGTAITIdfrfGGyOlhEbAnC2AJrjp8Wf
hrtSmLfmDtcPulsfEpTChHe8bn8siZWdIC+CaihGcHDKv63697k+c7KMo1QmxNgM
WGtqLRDSppGlqsCkNI6GKPwyC9itn/phOnOz53QabCitofMYomCrfZmFHVSklXyW
9zFyNq7jrXNFdwc3GB8Nx9rP7xt94cVSURPTcPEWilJ4pwYxb0JdeNzOfXgffJcn
to3++A6SethHHJwrIQh0WXaPFGogtsetJjKbfRK8WDsnSgYARvZ+vxGXEzLMTTSj
ot00fcPDoQlNd7fi+vlRU6F6mCusBGGJ4/Qfd+Ae6XxGjhJmvRwfM3lQobTECsLk
oFx0tVQqEJQ0eV0W87jxsjwlvfOoV9JcWwD6mGxN2vF7h/YbeOxfwlDBh5J7g2ax
3byKNQkQN2/DXQDjDxaQ4c2WqtMWf1xaTMiukfb78pXHIIEbrtsojQ+1WvfOZrTA
ad7LIXa60uAMXWhagopaGU0BQMsSA2qDSdVSy7Iif+u7zWinvAuIIJFLGEjUdV8d
/1WjI6FS2kHO7PD2XobLaHKsqOlSERzCdw+qfIBocjVjxhUV9lbcyJpClSrg5qSJ
D0Dt0LvFoSrNT7Vy7txJMF/37FDydD3k1YlUPM7p5u6P9SP/gnlsboXFCVy4Cg76
LS1eleGq9XQz8t3aYP0pNpIOSsIQ5piJc0fDx/lcnKBS+ydaiEKcxjrnRp0MfRFY
RQaL6IOrK2XJFKudZSabhXXEx2hKvi5CEGBtw6xg1/25TqAJLl8OacO+ogo3ckxS
ZhyGG2BjFuTmLbg7KSPiPWZhVW11Vb+OpYqJemhtQAk1wuvJvl8dc5Ox4MT2wfPB
Wpw7xIKevF95iwtEtbb0zOcfCjzvlsbt9tkACn55ExyegoIcufAd6E2wwW+dGSkL
DZqPcdjeP4UFSBpgDV7vvy696frcsvivNbqdDsVleMHf8bVx7P07wUocsW6ZueWM
6mBOH3+13MfJmH8jbTXtm5OLjJNuenWusZvuS6bUBsqT/wEjviYegzF0WjsaEUAs
E2+vn8ms4UUbapGEiv+AzARiIr4D1i3AC5lAbBZmPNH4AqtBGzUTnEl2n7/CRtyG
zSkG0zMaWIM4JoQCqZlvlVI1zszpw3eJFh//2qXKlIqXuQbgZC4enh5sZIXwYUa6
qZSHrRXYttu9Wip0QWncH9reVDYAvHTX+dFD5ImZU719BubTLjynzDJwlYzdGi1Z
8NDqqWCeCw8OxBcz8OplI6yvFrODgENuv4JhNYT1/ZeBxd5O0t7wMYx8AApsoYq0
dI8CyAWtEKK07XY1HKNgQZgSaITroZaa6w+nl9/7KXsGb06S3Obcof8hKkqTS68M
aN4jWok9ywU/Lm5jQ3SSCMYOGJyYpxr4WXiiE5XVkMlqM7aLaud0ABXUnVeZpZdR
7CHC7HsqzwRHQOwG2sX+5wvqS2MDKZR4h8HTxW8sb0qaiJt7dMEK5InmkANUIt0O
kncWhF0k51i4OFr2ixkHwlTlKucEb5/LaRo+yu2oeIF0lwzfHFz542wE5zyG5baZ
f6d3SRM2mi76lKsirY+ld3IxiUSke5gVbnYe06CIomoiFTJYEArwJTE5lKSCIrt3
locrQNpwLxdhejjJypl5Av6QU5zx0hWvFZ7ZOC+JW3/AS5b3MG5bElv3OAiq3aKo
ODZiCrU8N5VrVYviKgzlqMkx/fbF/SO/A0qezWJoTkcSD6YwdXAhV++DEwBRSm5Y
gLq44Mxk8YqEzt9n/ems6wcBd1AQePWc4ShRD5cmNXajyb0fScIwARG9I6TCt38s
3C70kCaQSFB43QcKrAe2T9uWMReIgfoZF5qFYI3J/h/PGsZC9E4oCsaCTqd6JJwN
dnZddr+X82q1W6IbQfQu5bz/EEBKaLwGuh7Yq9IMpmQv9E1yZBBrqag/FPuBgGio
Kysgfa1Inj02q14wkFw92moO+HbzFNkwNXj1lzvwHYMKoA+tosZECACMP0uXQi/B
0YHVkrzzLyIyMTlZG25QEQqaR3g8DQCX9Gl6Xmq1k+VOlLtXVqwewFd4ZWEwV3sF
k2UimV/jw5To0hJNLAHJ8qlgY0pG7M2k/hHPKekh/b3i7NewlWZPXPHxdO/IGlCY
fksUOZtRQExfXaoFbClPERt1ZGHP+lFTQCH/LoP5XdTdW8AF+zM064qI5ViuUSQk
a5Lt5u+CLJ3Bh0mHrWSlCbCCrXUq0bMiBgpfXNmU8MQKyN/3DNB6a21BGU7Y3ROQ
Jk3ZKG4Q+mkop+nyATbm/b3wncb3Vb2ElOcxjVmnPpapl4cOy8TX8jwRBZKwhvxU
Z+1MJ4fmmQW2s8EZjFbzfHuN4gSVNBV55uT/l5ntoDsKAMjTE81pNjFZvGwjJgVx
MgTnf94WziWYFtwWeVTnTtt/Ug12kt7II2o2Gf2N7LP5n4LcC/6a+bz87Dau3byy
S2jHnoYfpqAgE0nNSBUNWQn4zupFsyuJ5FuHUWJiIxB1pPoFi9WXc76BLU5osWaZ
LZF2iI8seK8YqicEkmFdd5PUMJMHbQVCgFKnjPCPEfg8nzDuNIMByLTdqH/xMPDQ
z82rxbIGKYZ7VAJVt8tzbqMvYtLMNLdxu/2MBSJeR988IVFT6u3gcc19q8v73GDx
i7q9BsaVlDj1ASAbYZ7q42qpArWzWBjaW1JwzcRPto42ITGrC6jJIuRi4p3+GxPd
lktaRGIHf9/SHaROnnveCCg/NRi9IlN8g2MvHAGX2qrHTJMwfJPiLuJks0zz2ESd
1ZKINicpqbaEKX2mnL7PNLjxsUHHfooLOzEYQnknzPAiSSoMhagBIIUMWSSmj0kH
jRFCaeNb4lDe700RVwZHKCN4gkHiuh8o513dHYr8sYy1gHHRciAiMlZwVC6gSsY8
ahll9fCjvyLKvw/62+1L7NfsoPLHPAbHK4FiO2FHFd8f/UyEbC+6KzJVK84f/Za+
6+nIMl5/oLztPPr/TU60gXjvwoawDthO1uOkTkqtU/3M4/FB6UBFD7W92VvyXSYl
+9r86EwNdHE7rW4Ml1e8IgeBJNi9Y3dG6QUR67piw1fLQnG/NiCIcxppU/W1Vtl9
22n0XHzrm2SlwLHEwKcqlxgSx58FzFrI6ZBTETQ/zKjHwMVrkNveOlBR4nsVXMBQ
r1+ez0912BbmFszJQsS+lXiAbycQVW90KKou0wqRHuJ7RtcMHGzDtXkhFk+Q55jq
/yIAkRs7aKNcJ19E8baF1rfexUd57s48Uy85CyQqBQENXKzxkEhYwhjUeYJ0+4+d
YcmfDlgQOFYzeI7C9YoerMwZNwXGzdzFL9PHUKoahMoX1nFc30pFYWX2ftHzZaum
P/zU5hpvDpa149SGNIsQIFyya3pBPSJJJJzlgPf7RMa1p3Fd3GP/XxeDQ+QSFIPS
lXgDT715DTSbw/lgebdFT+7JqipxYnlkD8AjFN/FJhV5BnqrDhTlfqCUHhmOhFdd
5wJg9T3Gw7AuI9cniam3w5dtwOops50iZlRAMktMdwn3KvSsxABx3uTlm4aaihDP
MGEpRiNnx1DM7tUFXQ25I9YArZg2nyrNYXYgqWveDnJoyElfb4n4yOLNzEWdzA83
BfLdBFNWQSFiMFm08dcXvapkFO0h7b4LT9Dy9dgXvh6B2MayUlUDmZzDude0aWN3
r8rVn9GmplyNuOcaD+VKe+CO6mD7iwH0mnwdSFXUjDKCheMh2+juq6CX10hZBVud
+xzP06LKM81UtlWUNRivsJzftVpp9ZqGR0ZXTHatY/8TN8V4Clt9/6opaoCfnxFX
R2BKECvpV+pLYhKh6JoxXQS5+rv6a80Gi0JG5o2HE+aEruoI4kGVopOQEtLPz5QZ
BVNj+JjfbhUFKaH5TED9WRmhVnMkPFiI+GQ9EJUKHbSTraelkpOy3GUCz6stKayT
nCZwP8WjQNw0KEhPGEVj7f42q21o7uMBL+g/LKAH9qyuG+dBWOpMB2jMDIKiEXwa
YRi2Z9Ju6x+F2D0o6zC7IJ0kBc+6jN2S4Hhb14xlal0iE45uful0MeoCBanHxy6c
NGNQiWb8cklAdKpJmYs6MT/tVwel1qWDs6AM1Qt12q/ZFtX3Eczt90yrC6s49x0Z
DSbDqCh+8mjOf9vMBsBuJ6q/ZiLQlPMURstWrJSagFKqyX6siKxQW8Fqcc1bEiKL
ZA0n9PwbGdtM8ayhbyxq3ciEDt5ZC7d489BjCDHPUdThmZ+dG9JHFARIsZrDTkGV
PTVExvxQ8/KfPpcZP97NbkcYRgKZSvynOwQsV6RmyZPWpMvdZm4zDD4hO6Fvxthi
73bqkxmphhi1Ut298vWjj3GfEC6ybnLuf2oSwWBEvX8IEPScvOWOhegzUXhKxwHm
k1hoC7wRw8HNcdOn/yjsLnG4hFAMijrSkVdGC3KVVpPYIzUq2CrMeyHcUwpededR
gO0dSlWYuDaLYXpYrfU/W14O/6E5rvmvLIEDtEwZX/DmEp/YXrsDE+3bfjGK+NaB
5DSyTwCRQVMuEIOmNskbpm3bSC21UUCgXfLlo516kZbjxo1vb35nNzezc3/IWMgd
dARxE3lz/zUBlxryJ3Vj4IJtHlhnS00YJdPjtHvicLRQmS8O34/t56g5hDlCT7Z0
3JgQFxnZufr+wrc1C6ZjmvBKXivTbK8rKVosyAx9QyWfjNzLIkRqV4U5UpIjlIC9
d9FPhxy+GAISaqbxYk+0MblR1MHafhI9MEV+THl+ARKtyQqrrbzmPaR8Syo03p9E
ao4auFaRbBH8jpwzyB1ACxOuWM0GtzagdJnqGa5m1PpfhtZspZL62aG+hb8GvpFk
6KMYolnB5el7rqwp4bbh5nGDs3xlwduVAcGW2gjTIizSzHPZ9i+W9Y/E/7UnCrEp
FPGejY3n5mO3Pfa3UHojJtKkxCYWnTE3n3PLZ42zbpqE0CVlOWOllHWaZpkRoZ9w
CSj5oFx7KzIzg/p9CmCvYVD4oVDBBkWxo5rjRVAxnpwkHbUVg75sPr7XP8hTy9WK
XCwPMCBfBcDO0Y4uy+mk50MEHN6vHHgQC8HYj2ZboiEMX39QVLTz/j6oQS1kzVlM
WZbDbJPVs4lsIcJZsSXsMAH1LyAAfiyad8TUtcrZjU57F2AV8gx2pSzhFOIXfLt7
Ywx63ZiqjrGAN35KiQ4fTGe4MxLbgA4teAYgEsmeRjSSj3NOrqA/Ex1msNeFB3no
dVmh+k/aUmQzxpgRizXqscJncsBUZG+FxD6niMSXmlXlIV6A0cSWelNALtZmEC3H
e+vJHVera41yCsv2AZ1oezRJbXvKAd8jJPgyj8mFmaEnyUotTfikxWUEZ3bvJEUp
GMx+QlFiIgvXoXnxdPZOIfJJlstputECfQvRevYeqe+cMRi57BGhm59mSeIqqgl7
oeqGU7O3Tbfo6VRebPsggWV9yu1MqvTKDFoK931fSosXLZU4Kazl6m4CMmoErKmJ
9mrdW4Y5VQMwgWvO5ofpXxfwwSoUTm8gfJ1Pi+v7rHfo6u6KBrApOPFcSjzmxaP0
MU4s8P1XbvApLIEmBJl0dGZ/JPZO8J3GxZz/t3Q9Z32qtXnz5P+BBEj97LJ2JaQ2
NB1T4a55gMO1i9BSHoGHXI+i6QUnLWSeN9Z2VjyAeqcIqOy+aRl77yhG/yIAraTf
+pbEG8mmirDHMlgHnM5HULfgHQtaUSH20x81AAcSZzUcUy08rYh8Alup8XbnkQym
7onGMK0tlnFGgjHDUfSgdQaifK1XjbBsGtIODm9/torsJdhVJxCNZ0FLguviOXNq
6sEbDQvOQgePzjUVR+kI6b7sbotffoJ8RcmflEPP2AV5UawPwS9MhpgLpGSRD4H8
xzdCGbgbNS6jadjfGxA0Kc1bVDbhdPR/JrdQDpFb4iuROQH6v82dbD6FKoHznOYH
V1zw5NulwKx7cqh+YhSnALrd0PwBlZfp8xUwpTc27TzGoUNz1juZ4CIotcuNCKdc
zIS7ZPru03pHXuzA6tLOW1nkwZHmzrNhSOuAGJvG9pa5jpRnprHz8bm0z+fOwtkK
JGApzIDpMNNqZk3RoA2Fa087i/6H+faaDPqMJjiJa0SH4js7qCqKNdYi1Ig/ZKDz
WGksB4y+f1S2h/67Z79/dM7N7jMI5lrjGa7cVvIGHkCcQTMAj6TSOLABGacZm8ud
YNJeqmYB0EB5oNNRu8HmX+sJ23q5q6kCVG2aeaQ27SsfkDPuTJZRxfvctDSMN2XB
BbmAk4k0Dri7nwQ9G2TogoyrB4+/duNwGpMQQcfcST9RzBFuJsRgfyaGd1iY55Qs
TYbLvp7WP/T257SZBVt0rWMqPdfH6aiK7LqMvLOu6uTRr2hRNjimF9daXvNS74Zz
uf17aC4YHkpY/KRLONwPje8ZSmkcwUx33XAVOkUvcA4b66YRMOjilKfIweb+ScnN
IlQFjeVx5j6548vi7MkwYpor6FPLhugDhI1VPK9jiTINllSVnm5DKD80zwYXlmnc
th/nwMi4WbNVPOnC/iD/lzg9P2YfiItU8G27kJCsntCMCa5y6PzzIL3L6IMBTWp0
nA7qjv665sE9SQGZa9lNGLWmvHhblugvMq8gszBUd2u4C8LmqjhrZF+DVqj8bh/L
sO1pWPu67PJzAz8joUOuuA2G78Wzz4XITIgddrks2bYSLhMen1/FaKcrsMO+xECW
MfNdkXSt+OXlEed+BfdcYPrwa6OOTVi5gmW2A7LwuhmDG9MePbPpCEkJKT6zHRuS
y1hq/ESGpKw045KsDsMjJZnLIGrBC0mpJt+2uuFWfZDfr2PZnIIdn8s8x2Sh5Tzh
XNCWrqYb8eLKyJLOVuXUUiskJdIBW3+rhPDfoSzV1sfbXpyGL13K/kWbz2xhIhga
LoU3IiUcCsKtRVxRZt6DkrGM63qZcl0fRdEsMhhHRgC6m/bnqrjtPtgxu4jKrR53
fuWeF/7dQ7RInA8QuCNvXoTZR4OY/6YKF1JMpN+fO9wXeV+6xNgwUo0plRv5Iu3U
WeI1SCqLsbSnow2VlwtV7d1bAvJ1yQ4ByL9RwBqNqi3f/Psi1vVEC0+jLRnfWopA
PA9Q48Y3MS24rtB1USh7qocXSQTLA+GLdf2otsTxDIpB07lNMdbZyasjezVMEipA
TOb9828hV2FgU1qLpiyDzzfr3Rtisp+1mxyZvE63SwXypALVpYJSfBFa1H0Btv01
b6w2n+smNaUV/P5vD+yhbYkcl/yVc1XSJ9oorcyuWN7zjt8oeciYydnPAN3X/1qh
FnHDWHiF7GAlP0nXL/B5swhVB5I5TyZF5656CpaNDHBJ0gFfopCer154LAAtPhOw
bhTI2QX/K960vhr1MT6cFnyJ9jfjs3Cb1ZTM/wIMb7eh/6G8MDHncwYmgyWwiVoV
cFbAnDAHBFLoJT1Sb8TubBn3NvYvyNILDdi0almPlNhewXG1/PcJ1tBfgpBp9z6p
hzH8rLZUNcC6UDc8PLMERsoQhZdkpx6A6jhAFPFxormryis9D56Tr82T353gpzUv
Qd6szZj7vQi0Zr7M9keCTl9Gerxj3QB5PaZ9ugcLGs/fXlX4jCAisbFID5NvW3BJ
iybnVEH2CHKzynuL2GFblxwlIZC1s9RlBYXjKNNWO+NpXCmATUYrqqcvhF8pPisE
9T7MGYF+/7V6OoIEjH7D5LIsY5OAAf+5/QA1SvZOGygjczrp/EXur3gUJHaZkOPb
Ab5UXT7242Gj34zGTwA/L6lgFvzf82PTWTmBAss/vWqGyl0xlGd/neIKXOOtyo5K
lItug8ANqkc+wwqgxyRpvuBJALAA9BJOlXHXhupYV37qpwkmKFC32xz7Fga85vwV
62/PBo8sjDf57HUDGawN9uXaJ5PzwXGRouX45PsMDdCP0rDAmcpuBghiNG1ZiaEU
PyNQWPohcDd81fG1vIkcX230zHhj5usggx2Nclcz+DnXJbtXsTufICsenHDLpFIf
fWRBNYClA9yywJ3DGIA8+BRpwLcPg8wirwB9FX6x02XseH/auLeCcKy5gKbVrlbi
KFxFIROITbu+ecP3T9cmJGE1/LEixhMe+RCm8wQotpw+KjMO36+flshfJXTU0mC0
aOAHirAppLiq+TdXFtIUuWPxnw67jY96AhXjmLF3wRrs6Dci2KzWCjulASAadPMa
452GyX9r87JsqQAcP4r/ssHJVLfaoA0jC66S1UUTJgla4jr+2vcfPWRwzMacH2S/
/7gM/rYbyHqR8ZDBYuAyZMOOKN0S1sfSjiUbH0V5NnE090UO+nJydAnsxwuJ0wBr
HRzZ5/QaXWOIHamsilGTFnl0CXaE2xuol5DvGWH03wVc8fAdObk7i2M+rCictbUs
XzFU74FxrCztw7mGqxT6yT/0609xbcELdlbK8XTAX7pINN/s2AR8PKevxNFQyN/w
DuQTyvB7qrDGU+sQOu+SOir2xelQKGK8Rm7vvjGAhfov2mDJ9CMHoHr+35EcC1cJ
vGShSu0PZw/g9YPGVwEbDkju61nwAxrWN6fir076mzah8zZc3nyQL8wC3XJQPP24
w9lLc08GyU2ib6k9sBWDf958guXN8Bi8ZULmjh594TMkqsg431DwiLv4EVYZDJDj
dMU3FiOgwESlEJ5ky5uvY5fVChvQIoSeZHpZ/JAYiRwn+kFL0AKMX3fBv+ZwytU6
h7bLZ0ft8Q7bN6TonmRfmAcJejbNI7GeVQIVzOnxD5cTr/luQgD+zrR4PpLUaH/4
/aDbpt4PINAfvZcC2vYZHaCbOQzAwytQ/VUGgoR0Fb/SMIphzQQlNj6MFCLZ9tL0
hf+NdvGIGfRKVbEEZpyZdOE+ibrQKy3voDUPCjMtvc1UUZzGqAPZPPxQ8usDavCm
+sgXanVVHsJm7OM5MJdDX0zsY4e4eG2vNn01xpYXcBQp1u7V6jfy9Z3RemXOGhoG
PVgk9GSN/YG3IayxHJLJjW2iEdslarnQZLYu20VkV3hyRyJq1lUKEQ+kyB+q6hdJ
/8yFFEP/FCqi5mY2aQtrxv43LuLBkzG3RoTxv1IpSRMS7wE+BOeAuTNFyUW/WwyQ
5oqdC/szdzdmEq5TuY8jpntxzn+8cu5lK+pqdORCgRUQhyM9d1PKAbVh1kjbVH7J
nuNXeNx7+M3gJY5o4+O2a6EvZqmOd+aTqqOsIK4sCoDzSgrEQG1S3kZbq/+NrNt9
uU2T3WKRkCJOG5JEqYR1sKcHn1LrqZFf0hwY4uydc9fbucxk/GmE6BMxMPDdaiuF
Y5apRad9CdiBeuo2Yfd04tCdSh5YKr0tWZMgatSn+qxpRs6nDiHo+RWaofj4bA82
U2XK4EHwWAlvTROsbLGGx0+TPZIXFPz6hxTWYmr9d6ARfQhUaHZTQBe7JjamolAA
0+diYODRZtQKdwTbvzu8GEYSeBQPujauIMQT/FoJRviC8/2ckyyyku1iD8RTACSI
amy7XtgdekZGaFf7UbYcwvxT5mHHxpDIuU166GyUrJ8VuvGZxqIYYFaLMst/JqRi
VGlCTFGqf+ifeeNrWohqYkYpOvp1O9d5fX8dApS0ZvB4HpqEUkuWp2Ok7yIgACRW
fTAEb2iWlNWLfBk5IKeXm3GOzm8akljZXhGg85SCP1KtwUtWmj0Be8LlGwY2dQiL
AN/K+lOpIOpXkrVkbNSQqMM4xo7CxWfgof11hlpx8VhjCQ9uf6zvjubYE+xCKWWv
dda4/ywkcia7JB9gkCg2K+XDKNe1/94y++4sFzRoZJkxobJcvFTftI1C0Uft6xL2
SGdqK/WIQtGT1u0RgJxub5TNDvdrTJ5K/EQtzSusl97nXx3Nn8XFmWHEALmFAL5C
mrAKUxulvhqNtFmbKkhe9VL6JajIqnkDjhgGmV81WxhqBO5xu3fKezI9gMVdOUe3
jtwbjIXWjQD90dZ7gPxb7b3JYxPGq1fhFB3sGsUMa4ZXMhjqznFYIFhhaaDEi8hC
7ozayCteZ3MkOgpQzX5k9FAxaVCGuhVJ9YuC8cH2+l7yvOn1oaJgbylk4Undpu2j
AQp8vMlj9jHEgKuSQw6Zv16BmlqqfIBuEDgjg0SX9fkKRXNWhNQNjIv/sIjeMYIf
6gSXbsubqAiD9Um/lO3iBKGoMV3gf4IBrWMtbzSwmz1kPkB+xmrqseVToMhKevKc
4DPeT6f95oVGvRUYO/iENEY61HFaPNRACAnKmgtHK+bceRumTDmLLnyKh+qevZ+k
DnDVH1zoACcf0fxQOtVFrKx4axsFYYmZnQZBUhf9EgfxK1eyqW+3cz1suKrkY0Nw
9j/0s7szms5dYWxJIJ9cdCwPv7oIzBmwXaEmFvsq2rUGvsc/gJhoL9qVaxkowEJ5
sFOxJhEBsnkowNtnzQyTTeMPnOoeZAC63S2dB1g1P1fCnHnRYLMlqOpWArlQiW5j
wRmmgg1zHk4ANQtxgUDD2U8ZdrziAJ4ZwYQXZMHdWmToXSkk5XvH0M/Pe66eKzzy
0LBOkrpludGMg1ljUEEHc6Pb6GgS1TmqKZQQTxwGBTeUclmiBhdfwKcvLwj81WbU
/Pwxcd5Oe1XvcmERBVr6REE8Q8/My/rMYaCN8b9SvJAXi5OJarmd97QjP+7p7GVf
pbrP9cm/c7Z9697ghpM/KgPAra4kHvhTZcUlEmjMsmFsWF9vKFERcmwkDycngBDo
ZNoQgIO/D/r/K0IDoj+ZtaUtQ/4Uz/MWoQWsFttpcMe6u3ijgQpdFZG+06jI/4p7
u/1VFl0F8JC96FVSy4Tuw7B51QKPvqEKyJis3X7S5X9l+tECuJJZ3oQLFouUjW5f
FE45ic8F9hfCNCRGUDGVIta+MGSPjMIFsZ3LKYLsbG+nMPLOFSFzZbnIwNRdnQnw
tVf+Eyc0UrBR/yxt2WWv584VRCAl3lsjKVeZ1Mn5+3XrButKmhPwAOnAf9pVIF/k
jHG47c0G+UscGIRttcRe/Df14oeT/uDdkrRQRE5EHfLl9fAKgC28Vcbv64ZudmOy
hbQqhpGzt+kGIxhSN8cxwXE6gAVN+0tJXXHDb1rNXtvSVD0CKrKIcuUd1ENFwx2b
Supt0GAYPMxFOhhiS+sAOmNL8MN1zPCtDqH5RiV5a6gUe1iLj9MvbRGE4jr4Na7h
U2zxV1cPKsM7xaXQo9BaT6fa2IgoAg5vAd/zukrPz4XCQC/Dn9o4QuOE30I9U0l7
iGnhiqmqTNielEfbJIC6SaUJUyRyKnmjVnywEBjGFJ2NwZEE/ZxCwGgCoUfP4UIB
bi/AD9hw0oCBslZE6K9mWvyFG53Ujyo2p8/tj0frIBKtis2CPWkFrLF6LsGYQfJh
VUnv08THSi3lpyrKLGSaIJ/g6ka0XKSY1vZkAZl1QgGEw5W2bQdWKq9toj0QB32v
XexjQXOUmd2AiP0eGmzly0+OP6g0KlI1B42IYE581NL88xGVemXh4ot9zV84Ugrp
866BrgXWCjZiKaZWGmTyU80snIFKUmlRnMuGvPbHqhgbdsdnNcFO1RFZ3GPCzjuQ
pAbHJkQnzrXNK0yAHnFvYLHvPVapiGJl0mr4yL5IS2LyPqc3G1sDBrn8Hu3n55m+
N7LjumO4KFafmu/E643ZL9piIN2VqFE3LPBgqNhJznW71d7D1GgBbPJG4H8TwL7T
fUxv5v7AWULmCtlqD/Hk4CGES2wZ8e37x8WzBB7knZcu4jXqVRlKSxQFt2+KhSGA
4nC6amy1B8YNYBO1ALGcSxZqldX/G4p/jyIINmrq8sWfVz38CBaXmC9nsXa7Qi6z
HBBSuNi/AvGCiqZGnPtYEai1uoPb0Ykem9JYbnyknSVisYRCqlGgC/zNIr+IlQqA
fo+mpNFF6ym4NYDEu1iGln8bwx44QYWx67vaaMkMcV2JPnJVvtn3vBnJl6LSAdO6
merLshDPRA30QGj8IIrgfxyqMPEF+5iylQsQ6xOCYkRhIaLyEKV+pXWgz0HIYuR2
BPRwfu/qI73Zqxy+j7gVVK8+MNbGgQzY9mL6Yhi+3dAxQmd/3r/0wux85YXx0iYi
ahYLlFqMhHbIP8VT4G+4PPSSIaNLQWQVlgoklhbb2iIG8OL/ymyiLrtxY5D6CZK2
g2qP4y34g+NPOQAjWp44sAsZXQFwFa/RkW/92HEUXizz/mfMzL4P54aBogKSV9u0
/XQ29uMBCOfLsGVLBNZhAPnwb69z+WobH7oHKEOeOq2v1AZOrb1zfXTSRXHBOmTT
8BNrDklQ1ZiIS3KE3nlZAp13T6iyWku+lOxXCIDr8IYdM5Rk4gNuqjM5p+mrOWJ9
2T+ujEmHyEaQrh90do7OzHbW6nb/t7BucwGPu6UEdK5vf+ADBU3Yn4w8Q9bhvvAd
8pPfqoUHynshuloLEwbnhNiDvdmZVVlYEYQQXmnkoqOirjoKjcN52D+ypiAOychY
+uyKuDBPlkeBSmeXTP5D1eF05BBn+hCruTRGp8sWDRv7Xxyj2Uxb7imv0a622qGu
vOCbSfLjvZxp7vs09pSNeVMiC2TnLFp3XTARP/J0CYpU0XCvAMQvz1tupw13GbNw
GXrl0ibPDZ2EPQ5WWzdZ/ibvMKZx6aN3mlZYCaUz6C34aAPNsMJD5q7DA5xArItN
yKrHZet7QE4LSmfCaXxvnMC1GArWjGlRGmVa3kLWMBmNRpgjmMoKhHU+69FxujzZ
SsJRXCQQg13Q+REc6bxwIwFZWeplkgbfZCDzxoQcRP3nrNWPccNSfZQAucj5k4uS
iLDH79ffWdR74hxoj1W5NF0ezp/7j9fouY8JMMzrAl3vSgyz8L/4GU6NCXl3+Ov7
7D+zxxGPneScJ6RMyybAVKuOGDdnA+RtRLQCKUHHT9siOeaelQFCizUxapKyw0yt
ABz8e/cZShByPOrQHIS0rfuXh/qkkd/nZAAanb3SZaDCFQMR7oLIAKYyLlBk0bV5
RV2jgYtxvX4WAJPr8wyWnavr3Jk7NcG29HOnh6r5rSSVWBGR5VTv9Ft/sv3svvjB
ttCikRs673k146yFbiPEDQ/Z4qRLmeN91HYW8R4YLA1ssuW7pb/B9hA661D3IOKp
aiyds+hZ4OS3z9X7ijFAAYTA9mAqpZV4KskPSUmTSMT0IvaoeMjSh+SK0QIT8P5l
2NpuT3I+mX/M4wQC1ponJTJ1UJKcUZR794NiVNZVO+bfFTnBjAXvN1aagKL5AFbZ
EtBPqEmMfc559xB4IhbRFiRo8ueo/09zLI5akd//kRTayUP/iPLHv0/1FmLL5jT3
p1MoWGYLVgYz8rkrZ6BTOxSedjk/KKQ0YJZUQ8Y/xTnUfQfApZNw66Aqm/jkSRdc
2f4MV0GyP+Wy6qs8C8Q/7UhBi6h5izxWIOQteHUpPaQrOTZECTp5Qq8BdUC0CJoi
uzxaDdQu1jySJjfbl5+atej34CZ5IYV3l9qURXicjQ2rvifeAP+lp8fi2SIHpnLq
6CA3TzJfwT2Zj8WMoy2N+eEu63iu2lgLySIHCtglGU5QG9u/Mwvgc3sMO+YIGoYy
TXid3lYhmIan+Lm+d0yvbuZuPsHYzleqcAfp6BZ7mtbRlzcPjz3FH0kd1WLRXzvL
pj7yQB01ayTXH944nXT9/rY18/Ty7enIk+KNDGqwhANBZvy/Gaigep73yfZZXRB8
AA7S0Bn16Ne3w6sTQ4esqUp7Gw7kP0WD4AtjxY0fwMgcKYp4041w4F9aklVgWQwW
Jq3nll5Nb3l8qsVme6tI2vewl2JNCB56HOnL06P0HKH92MNWrCOdLQgyqnSx0LGE
z88vXc/IuEMrwbB1Q1BcKvXobJYQ0B/b5oAK5tWsaO7u3an9JulCjcerxCuUSjxG
zj52N0XyvMHPp4+BImA6VygXQJUgCUjMGhNmjijxG6uAi0mOjqoygOEZcohCmwQC
wsJsib0fCkT98K2zRJosCDiIbVL5KcZEAgtSx5c3WD8HlOMoprhRFxGk/pPYqSfM
HD43uGCVYyLIhEZ0S2QU3aNCp85CPS+9OpxNTLDGNk6MtP8rOKe3E3qiZmN04v5E
Rwu6+l9qutMdlJfhmoRR7Y6MGgsfPQx01niIJwOGKayDQvoAl33N4jD8mwLAh5lT
+ih4OXz9mcpFcF6kTNgTDOvsZ+Efk/JIKbeVZ5SPWhatLh4QMFxwJH7hFr4VfA8f
+OBYYsu28ht6+qSKAzF+FpOMX5zMn7Q2qay8Jp72f/G3P9hP4R+6OXdHPfDG6au+
THicHhDhKeFMcIN6vIYCHaGshVnJmeMX99Bu69ptRpB5F8MsvNiV9pXUcbCV7jZa
1o1bku8rKGeAzObo72/86VvJ+mUj0WceI+xEooCO1kHdwqqef7YkhhTto/VuCFtN
9Y1NRvzn/iowXWO5nQv8WwBKzogEXWMIQMhLLTf9sb3ONHWHIqRdDVVKKhmuovrD
5dl6it4MiSXU9B0bTE7wOFwquCogZijQ0gW/YVrVchgA0wKqLFXfVjNBQsInTKUe
N9eEITuEr8x+yTFlRiz9o0UsC8wtFp/TOsT1tOJpsotZoy6DU6N2Q3RMRh850IuI
POiIZQWTbOkFXBP8S2s4YRhJKhPMQRGdapCZsWn2i+GHHeFr8gJJ+zPil6LTP378
CLVtzggOZJEcGuZBdOI10WfDAze/NOamiru0oTiIOyxj20oqGUK4YDXBo11FNv6A
ioy1XcGgosDuYVjrU6jb4oorpPV3GjNgRDLrX1ezY4wkoDhgA5IxaNTIlx3wkXYL
38D64oeVbL6Dea/E2ugoVzjJmJnSpUjKvEtI+ZryTHWmP1J9sWye/OQ7X32egUJo
bNrhgkpgsLkpxniODgUlwq0ffL17h/UIEgp9onNHl7Ph1c8guRSkxhEYMuEsi7ys
McMav6r9yNYldCHHwaXZutlWf2IhYKDF1HqOsKQfsCHgntlg62aQQvRHMP7np+62
crEgj3qQnjUkkwmbZrzhlN7X9h2AHsrMzJjT8U9LNUm42opz600bU96g/COlWTRB
/JFBME7RVv8GbWCzyhvnqp61FJ+RkEouCjsvmnvmoC4wdHkqZWrp/K43UavaM8yH
rimY9bAW7eBsPGnI1iUETf25ruoExlEOpmF0BSCODsycDx1LjOxwd1BRpHgbXdhx
bBP3/AfMoJkWBXnglk6hiajTI3ZRfbFBrzJqxQ9BntIVHoNUUHfSo5/KekC3sUoC
GFc4biYkw+B2EAI2KHE706WRAtqHIFbSa5hZuPS+PGSAhUZ9WkLJM7gNq/pDPY+z
K2zpr/vRJD6TN1BOoAdBWAf/9trmtxiDN19qeqisFfjgwXFHV1A432KsESbGOyt4
HZ91D15gGBt/3rZajSs8cl2rU1iuHdSWdvlpkuqnmFcE/VzCdl1BD6mPXpw1xBR7
x1qbWjtVyeVpLkvw0YrEMLKTcccCkx0CKi5K5V312kLqt/DXa01656ZjRU45LWQP
1G3y69w8wA6PhiuyoYLcQLzUlZKk8rp82QDqpMegNzbSBifQWyzEqnM323QCcdhC
yiLTAHXfK8lwEXacsS9NKqXrsUVoO+Smjb1cBnPuVfggIQ2v2evBeAfVfNI4mBbZ
TOEkoeK+sVeHojgrbFqMFdISdkPU5Bxu/s06cdgSpUuZBabmyxg8Tk41Y5feOSMX
i8d8N4pqk1TAzo2F8RBLuiodaV9TqrG8Kc8VbwT9QXsMgYJ3qBYu4+wbRoZ7d95N
fheeWnF54IgkGc6jM/cdaWj7TXu5PfxtKzIBqL566+Ds0+noiMC8cNYXwWPBDDeI
Hd2VvGPIvruouErpdc32868tCFpa8g8SNf48JTWeyGsZf7HOVlrMOO5Vx8s6wsU9
x9Sgye1rJFxdn7qcWjdLfESc6NX5DbRU6lE5px+onRMDA7CY6i77ghJuYj6cb+gg
7EYH2IcH9UA7aSFMbYnyNLSv0zD2c4JFvc8p9nBfoBIBWiMHY+qheFgdyfFfzft0
BPoYK3gZF/+NtMcGg7MQBvrhHv3SH10AajPE+W4cStHl2LSeclXdhHGw0/5YShpy
C9GOjot11iqY1xE8ehD/8uoOqEKmPUYSUJvjj2CB8vqjrrIO2Fqtjoao1kdQx3AJ
22S2UV1/OEjuanJ4KOt+un1C98Q2IatFhBjnTQTy4Y2zoy/czGiJriXffAdUUt0g
Jpny6YPN33o4jguj9qEQ+Nq2EOFmzYUnCgHG5taeF97oNlUBlO7ZqBBJecW/yXuK
EWj4dKYvwzP+gPUZqXq4KagX5GRODZs3Ptt13eAzuafNYz5W3n1dtzHpiazvOYr/
WUOsVS42AsJCmnZlvK4fGP9gi9jgpUrCoOU3hKPjOQsebfRB0wESjUmD2VIP7t45
df2yGODjW1WoZDN89CRIazwUIU+5R8x9aLfmdjIbofhPfy/srRZXGAHJY1hiTkRM
m1Sl+nmXu7m7vGfcLANHoQCVRwQ6F/bOhdTFmHzfLLnmMIUn/FkNysPiFIInXOzm
c8nCS9pWCF4eMeDL9I4106QOQD35jlO1SGNuZIG4Dj+gSl7I9CGxBl4G+u2w7QbF
UrwaWC4SGvv1HdDqFdbXnTpAuEEb5G5fdGJX90s4OFdYUIlB4lKWsmMuu2zD35In
/b/TqUHHfHRt7hdLEdfPQRBYxlyq7VEUhAgxeI3d3LMY+NNZQOXJ91IJCfbWkK6U
uxdwo1KDoF+NFOTsxjfbWTYbCWJmbc+gAqAMhncQLQDI4yxeP82t7pYbFQOtf2Pu
Y0BScApI0Dfayd3fGnhB35/l4xT0WFSjfpY8JGN2QPBejto+4koqV4WcsgIC+zul
NdruKxrDkmTHaPgg5n+zvAgAGHnhTd2F8FN/fhb3VSd6pF68J6PF8NYnMTPIEPXd
UuGcpxJjv1BF8izyL3RFr4/dIPkTMlrEIdxU3gSniPx6lUoVKjy5v7n07bQcSQ0D
2b0IexCmbk7irrikmjE6EakXKSbBWEaC3nXJsQ79Lqg5zwPqxV1/DO15Y9whZSq4
10Rgj4QMO15rDF3+JsKu+raiNA/8VW80xyOmkTdOQ5cPzSYRCxe6NNwX1OXwrQfB
5LTOs+cy2aKZ2OfEJBFBtbDaL70gCDTnPg+rKoQgIKkYc9QhrOmpbRBS6fqA6G72
/2bOuq1Pn7T+wWic2rlpZt6svPANYkGQrlOtEngESreeKPjvzsY+cUslcz8CW60c
0yvDPxw7Q9/FnDONAiwSd6pZ+Sy0omSR5EtQWYyRfrwHChdGurq+MuE5ji2H3d6k
LD/hZt4KrCfL+kVCrGXvw3I4zbxxaLX+d4MlJtjc/URCFJi73DPrXPasFQXWyui6
evpdse/wrf5cjm79x6H9U6JoVWxzLuWmJQIBmWpFZOUzDrAIv/IBRt0JEZ3lgqT+
xvEejE7rdrZz9Bl2MMIKlRK2gtgyQOnpvObTkh/kE+26PQWURVY6VBkcwGCLAHTU
uShtIGvhjmoArcBG4+Bh4sqZJQSbZAkiHBG+UkUmBdQwQaTiJ5ORWHeb4MTlgxlg
ODL1igqu8gCRuvSD8B30RHm3o4uyTWlNBJSC0c0M0MzgSITJFo+8lwmTZVK7iIku
lJKld7/fIClF7YTy/4YfLXMer7JWwFi/eWSaUsDFBm/L/v0cL+wJ4XNMtQ4w2zPU
VhhHpjC4IHcctPXm4JQ8cRZIkwNi+HeZPg3XcqYlQRbwJn3BDlNr2HJAGc/CFssI
sw4SJNKbEdLxKsmHDJVjrnEOHJHeSKYd7VNhKg1wKkPg5MHcoqh2oS9pz6hWiXRD
2sZ3D87i59MX+pWMgmSS8idW7TGbQFiRp5AfHRBBcmxLSLWEhPhkRXhFJyPpaZBu
Tj3aZWOTL6UO99D7Np3qazJTcvr0S4bRh2T1Zo3T0ZYjCHESp9xRcxT89Q2Oz/xr
BeaoEHUd/Cm5DYJtyZp8r73MX2PLvAVJC5wa6vxO3BGzgmcFUNnWfrXTUqACxvOZ
MrvVoeg/pIcjca/V8n3emNT2KXCBYWe5aXLw7FF8EQ9Nia9Zb5tTYtQK1djVFtzf
7uc1adrE38ymV+tlW+8J6RSzBEyhYeUO4hK4Twkc8Sq/pHeyEOCEDg2W7Rv1xkBR
nR14GwGBDRHOTEYhjpRCyx0XVO3AGB9gFyghX8yK4gtzvC/Cv5r3a43mfCXB+ph8
udccdjsjOIFfPhjQFyjwMT9/KjF2JsA5e+xOA711wDWnAGUdUAX8NOJoCUuTqi1G
mdpdlgZ/AcWTpjqKwUiSIrEiAOTTteduycBwsHAL/wyysvOULkem5SNx49Y2CDY3
qDtNsIBRDGqEhumaCN9Trb58QwdBVf+DXKp2AfcaW5WAyZgt+GaDH5LqmZT/RfNA
mtD8q+YVnqx7MRjuMzqBKheHCdeVzxFHWu4nj/soSgrVTos0gOmTM06BMpECY68Y
KKIklQK3Wkno4My6ds9yt1QpOt95vm/XrImnOPBzP6g+4/KO3c4vdG6teXII58bm
jJIbhliGYJRGznfP6m0o02N8tVgBrpEL3yci1gTfoKnV9VHW+6JhJsN/rtt+JAnM
rxKeHPmsZo/FdIqMjFqJFMx9CTu+8hvG9v9sARrQMMOudF+0oOcApXXWM4mKNlgQ
YCavsI7EVDi0sdJ+/PEGVeHJzIDQD+uc7w9bkYejDBJMz0+onqWogE0lffZ626Rd
Vw9T+hGGb1ZJ82Xc/ULwstjzJCq5IgInRalws+PfPZujutmOwjufm6EzEJvdEAgm
kcG19UdqF+jEbkIPmyJeb3yiyOA4E3MN/OMGRqRgmfCXbEOh3X3+odiffUlgue0E
1CJ7lwReBuEnPbCDz/7SWdXK+bQhy8Voh94u9smkVL5O4IrOhDoDYekPCEzHx84B
hay7NErySGhuoFvUwu7K1R8qDa/CAVAfTcZ68WxBwTytvF/uS/Ptx1YP9ccJikJS
s/7VhLJhFtzG/Osouxtsb5YchRRLkd5b10d8LkD7effnTm95EzdQ0rp0skYTcPp0
XQBKdCl4EMwobyEzeyIWaWLpRGRrDXIZnS6NaIIMj1lbHUC+2Zwgbj6vS9EZMTer
a1iMlchJIWu4tSHUnoB/SxAopuh59UvI0goYC5OjofMnJv6KtoPORrM2czDxPS1S
74D+PuHYA7UztniRkDBwxOBOnCt9ygXwLhh1sD5a6e1A/q0Pqqbz5WVJJHyfP3MW
EDWxoZxOUOhyJ2eEOSHyMkVVv4yS725/UHgZDcqyBPLnjDwe51NSf1aQB4pdEV5J
kkCq3Xu5J2NymMszgMr3LWJiYm4KwbrEVrwIjsGgWIdktuoxG37EDGcCBMKg7F4i
HflZ2ToKbTTq8qScNBBqQ2mVlsonSIRMc+B0IwH7/NnjLrsvbid4feliXu9a+cmg
DYv4gX6qOuECgkZQutdnb59svkOxZzXpYVoI58WZA95pz+2t83sRD92nnr43bmD5
8Hu+MQV0W1bv1WZm4be3uvNXR8sF6aUGUVXGI8qAcgDN+JQ3gGH/ix2YvqXoyrIZ
9CYBUJhj63ePLkA1lLplGN6in0q4Cmfa4OrlkYUYPGe5Lhx12/zSy7sglUSaYRdi
bcEK8JFNZNUcNgZ50xv4kpeo2zwK0C8SwEAqR+35tKL7jPZl43vbGNkNwPhkSdRe
WSpXgNCy6p+7jP372aKI7CM3CBRnV2v4vMx8N4q1L3jvdkm1iwdRQmciI9H8cev7
7mkKPfmT2BBTHfw0CTYKFIF1xUDl+iGspF3Sh/e7XIEc8PWt0P8iy18m4srMqKBO
BeYNg4d7KF+Ds8FXFTFfq2OIHx9CdcZAhFgcjgkqS9SYr2LaflnPBHAT92+8KnE5
r5FGOgjjstTcyaBWvDgiWEJp3tr9bWLXapnNeBF90hfwTUb6Z7OqTX4Lkb9NwtFd
7Br6s1sNKZopm4lV0t5BTPVn/15v+aWk96voj/RncBLe2M2ii+P/NPTdFXvnysvi
p5xgz4LaFGZv723e2Sn+nav+faL9JfpsOsh6XfgfRmaszOy1hbmBlaJmSZUteIT8
v5sxj+QuANVAi1NefJuBOxJTCfkzLzaw6f3RWYu64zDnY1oE4gaDS5BUpayBg+r6
KyM49Sc6BdymO8UKh4axm1Z2yyJg4MRVdC6T6VsYegEj1xktBFgdxU7gpwytyUGi
jURoApQGfZtBkBYqRFyyGlYSzR021BuakjIO20ZhgSY9eG5JIRy+ygTrLtGLuUnB
CdRCqwSxwUroOdOe0hLsVcTwXdFT2UOEjrxOzUzSZEEfM8oGwD6AOtJJKLWj44QF
jivw3K2If9BB1BiX4vkHkfADSerwHoXnOy1vH4WtIJL5nq5fDgvB/iholwYC8jgk
vb0BoMembUeGpEtPzg/93JRPwV0S/xssV4TTjDlRDSEJGjEgIqjnNE8sUGy6K4Az
CnfvJtka9HA8pNqtNCfmD809W8ZsCyS0i5jHf6ljyay+byKCKjznblQFcHDO3Z1v
yIOe0TmdLFG5cLmhvQmEK5Cj+OS0u8u9C8M5/F9J0scdL6IJtQOw+aj9jxYTNnIP
6ytDDySl0dzEW4cGwZXMQ+TTzNopJ+geCLvGqrEvu2S3dsCs9b87IOw3hwsmDkyc
EYeW90QOO+qZOwHbnT7EwLdDY/hADwPDPL6nJAetljoU/4QKVqVOR/4Qbm/Cb8nw
TmvczxSEk8yRKiytqSIjtTodSlyvVeW4CKIFfbDopUO0HXl0Ep26nkUtHrBkLcPt
8slhaJe4rfhO21HKC7iKdwmT7wyC+F3x2cFYP9lIcYCH7BbBrncg0FOdVIWm9jFd
twlLtrXaSy1x+/g7V8zH597oLvnt6a1amGziwEs7a29BFxOQsGjiZA9Yz5w1oRXE
XlPL+SOaSB7sHwFfiVCfgia85jrCrvtrA5fAUa29Y9a2mB4qUMLSsO7Qc/Wjg9aS
YcikHQqq2Vm1jYs0Oj31u0mExixViLuBl3eXRVPOToH6ZsXCc6hIeI4ehyTbTqOg
UABezoAPVwaLzh/w2NHgrfV2CuKLz+lUg61y9MaXyC5V8TVU2cTj4u9eCTi5opSt
AopfdfEQck0gIo5Y9aLUna+xUQVPACaoluq7Ivi5qD8rXbj5QibZpwW0qaIlygdq
ZV1CsYvzqdScnHvPcubIBXNw5UOTPXvkveWryWFEYT/P9+ZBXY10MzkOFmJchPdH
1fjKQX8HZExU+OcBUVWhxuGkKhhihk/GFUPyhVq49R1BzUJha6T9DWY/io1KDMVu
h5FVCi/JV5h5SnWLi1ndEoqLDoGPA/hdOhONaSAv7TgUSrOgpxn3/6QOmMxGcZZ6
uDtDu2MmpyZK/NLriKBOWh4YlN/Yzo1K7lp6tfvfu3mmIB0//n0bYJn3BlLlhwXu
LNntLUyJKmJRx8lsKpb7Jg5e11uL/87jQ/B5gN2S80zCoxZB8FuE/E/Sm0XvZj1E
Kwp1RR73BUtuh69WnFFo1Nu0YMvkc7T5eAyCsknyCTQoJBZO+2y9cx8XIuQVU8eq
2JKvVEz0uTnccG3V53rVY7kcaz3/RNJNHo8Eb2T7INwlrZlw8dqI+u1d5esoip3e
9F4UxWR+lv8lVIUdGCpfXDePTx1/Wp7k1qv3db6gMkbjlfowHeGyDNuPoZGcy+5S
jW0F7T2IFIuom4DrSHSGRwd/3xAbCedVMnBKIVr8Eu71VqSST3Z3UuNZ680g9RRT
tRMHCd8rnahNhpR6xzGcUUIETs900jctLRr3gdr3XmGOk2t2RRkas3dfK/MXfCiA
5lwi2vKAoNeNE4Co29lcjBTFqrr0O6V22ykHERN9vBiUX4seu7UkInKWWQM94JCY
SiXPT0tu59Mc66gmuN2PntnnZvLzMxrV0QV3yZpCNGVXJNG1DLKVg/GJsYlXu8E9
Ll9qLESjlV4NrT/+B2X6/HW4LtpN7yc0VSlOM8Wz6BGE+Qh8+MJRpmciKP4IZBOo
ceKwFtKxzWESOC8LM/0Cpwvu487jTeE/02Vxnd0ARzWHxHKWm0Fq9gtv1IqliekC
AfcZyNnG4AYkqXv+pVBP1URrI8MeuWIJ7Gs3JQZOzZEN2aFbkvIbJbDg/CiRj82k
pjijh1zjT2xQI53l+GH1l18gFz+6cQYDPrYS4GXjhzPVgsHLtuUOaEFdo4cUE9+C
LBORsYloq+O6cxVB3nPmyhkub5/Ul8REo9nUYY7rgx/qWxVxmPN1SOGb1UAPWffs
N+aqFqytAIvSvNsWGEnnm44UmoDNod/hzqlzv4jRuRcEoZT5EOkHBgO5M05dAojs
n+twLW+PMsRq0tnluuMNHRWSw6tO6OiYwVHrluibyts+CupRAvdiSyLIRKGaMNeA
6FV+g4ftWvWlSl/70KbV6fATH8dKaykOnYhR4vq5WmTZ8wu8DzDw3pxACYnAN4ze
8Ucp15LV9ALRvtLPL/d7wvT4HjSoREf9u0gICuoGtaaBJiQS7AGC2m5tWIlms0XV
M/Vot9cYpkHSGqW+igcjbW6IQ7TtMg72bm8k7hsskcdb/NGYToIiSwtO8JA155xZ
TKsU3/8yl3acBJ5yiFe6Ss+C0teXHmOse08kBxIJqbFW6b4MnLxaegu5kL8uzVcO
01Y+yLi+oAIagO907s52YwLa2Y0eF/I1TmC83H1ogbibSiqFla8T/cte8jKdOg0+
IKQ3UKDoQZJF6U9lLeXoAqL36HlNu1n8WpvNq7EITsfJ20XbsJOXIsLXMpO9mYbL
yR5Mdn4hNfCrBwhPoLBQ8yj1GM0S8NAku+ycdvaxOuLuIWTl1rlZZgcF7zjJVt3b
0pO5ZsCldRIVgsNeVmMY9f43eI+DD89VdA6oV8JQZCG0N7sZ0487UqqAKW5aOBY2
4KgpnmOld3K7/pT0gjEdhRIEVZ3sG36kmHyhUBffUgU98fK7YckTvQ01sj52o0/b
geF0pdPHUXhxbUTFVw6uMrTr8tCG5RmKqVaMb83Upcm8Xwhuu8+9zUOWcXQlrFZO
83SJqQFxqcZ56BRZVJhqP6LNccEztpZt0A5l+XmBSheFr5IkJXQijVKCjz/ELP3i
Nm8fFGyOIRVCOrV4ScaPwR+14zDhg5fxnVWxAG0/QaPjNizSFdJTG64bN89gkJDW
A/T1MgmwUTVPe9bglU7y3lni74zpFqMWryWOBP/agwv7ndUnzz6eiEdoFonBRX/i
W3XGrx5M33c2spM6lIViA+zKOLzcBWOItItXG35A9ZxDitaDpeh7YRNwamQyVGX2
NUqX7CcuNYNrGNB4gFP6pz2KP/WWjK+pGCvCDPHuu1bkqNE11xjB4gu0Z6hZHLZN
w7wpF+9aHVsNSw6oJf+RoBEGJJ7ah3TZ1oe9WI1jxFrZZYd2CpczmHoX26qMbsWW
HTiDX+vUOJLDh17r+EDuJ21KWNKW6HvAooQR3rarVZSHB36UN3yWdpdpqyWh9fZ7
eKPq8Z3S7Yh7iq9ztspP6jZbUYswfX0Kh4y6EGNpcWMomL63FcWjeLZU21N0+Ki5
QAPPYQ4MtrT5eoI3r1hdzoVinS4BT4kkbOVCFdjI8KM+/Gzb1DTo/un7Yvyv6M+f
S67c/rqhyf4rDWvxgUT3Uo13YyI82c8Eh6uL2Q6j3CPrTWzvBQi1ln22wcLolV+8
ierYydZUjr/ijiFhnH3TMyQz3iYaA7cbyvhRnruvYhxXAHO4e8MmWVH9lJ8OkvPe
rwcBdtZ4vxZiwJ3ntydT3ChJ2Pl9QHMFMn/fBf57yzbV0CjYNemWvCpzVcrneyDk
jDlukTnz9fk3bR5GvnDqslkfuGXWtpBIBj0yK8odrCGvpB0qLy/jTj+h6CqNPOi/
uTeYHGxVPBNVs4/azegumTySml6GnYZjt5IAjK58exQeYo2AGeFnHQc6HdheXRGk
YunZXRSDqXu7IRSMY+GtA3dI0Ie+hOTCLD9rebz37WvsU1Pm6lTSRJsRmArc3AHL
/NPl9d4hOptpytmEcm/fE4wyfxF0nZPJ5PO6N6cZRB9VUegDuV690XawZjNvwCeM
Pdxy8zqD1xdpKK6a5DBopi5KllJLWawjG3843VMTlgaZPp2ES+4OrwdYid3vUWED
cHWtA58bHMm1mTDT9KLaRGSG412zUIpYRxhmUzCU1zQEOzp+39Td6JQjuNL5KsFf
CKs67s0v1cpwyDQCChtCuAzK9YoVy0fUFbZnNDvIvs6he0Au7TqlXG2/57pHD8R/
ks0Ekbg7iYZZXSTcFdkGIiurpz4Q9PcdSTA5cA3ZSkQVj4DtOU8MhkWjBOGcUIB7
ZPsmLft0KK/cTo4abSN68ZTxsiGlHflPby+/wPEXvTc0OOC/n5UzzqpunfMte1PF
ARnf90+PqGt7zmBtUq4yfLvs9zawdX8mSoVkQ4RYQxu6Hc8NHErzJ+kskCNnNFt6
nJ2IzjkulcOehYA2aXJBp77sg/ra0XaiYmZL2F9ZeUdOiAQcoPPLGWL+ZMYoo7HD
jCThJGZn1ktSKm8U31rxtyFbv+C73+wFVAjor37TY1i5OfJ2lEem0xnDJ4Q72o3d
GXgeUt5tAMCPvz5Q5rLDgghekBnTS33kZL3dr34pGIov6q27iPQUxDEpx+LzwZmy
7XkD4DG3aghYYTy0dz9B+qQkkYi9HCOkRjM0c3Jb5QGkiL729AZKIF6IQ+qmj8or
0y3AbEKwCAfNKEnbba7d1ug9xNV2h7sXg0vemAe41mcvJLeEWoODcDH4lu6eM0he
sEPypbYeHPV64CcxY9keUFi2L4V80F7HsS6TfE0uvEccUnEUii3YQYSo1HzBsfgd
o1Xemq2DodqDWYNExMFxl/MdF78CgKHQX35rLMUol9WC7BFsXUD7sd+BRzVhbKag
kb2RmjwN2qVwT87Hwukj7pqK4p91NdltTsJi9VeEYlAZJQlgWRVqpAhA/1tpB1Ww
/T5O8s7f5YyZSw4PTSoymmekzovbnZ635E9QfSeIC33DMtG35Q9UmsQwVP5DS1Or
FYXGQtjzxIxHwlw7y6IsTioFbvrd1w+CR0qrpR4pj2jhEwIfgAJQJmH6TavObpKm
VBS38RWoQuwb3j2O4Jw/YtgVkTq2+Du1WhIadf0PeTWAwTk5pegYuXJHDOsUYhMk
Z4G8mrFahG+YoQw8sH3kf3uT5C3VtIqK5RQl1WQfz64Aigt886OSEqNaN4qSC/gt
Q0Y0Jv3zFA2icnWTvZuvV/8zuAWfvhvuU4Wl2VxHGdO1NZx/wkeKKAbuu3Moimke
BoKuscf3/nn3T65dGiluVXOIr+XcLJsXOXA1NSX0vqyB3X8TXtjf1S3S85Iomyj3
XiWxFktn+4tWXKqf79hRM2fsaQVZDOt5dGrgb03atjYcVbQOiEExQXyY0ZbpTJ3x
wlQzgtHHA8u7ybkCVqsHh2XdVSzQpa4WdEA4NUIV4sMdxUEvI/igTf4CbeQ7NF3R
eYbrlAWRfOXR72odWEX420dQdXHHO0wjtseTn0IRYUfP76VnCS/q0dH/XGXRNznd
xcy8x+cU4SAUdgzvbuvusLFkiUCIphax8bMWxwxXfAdHerUnJDIBu0/A/+qv6Ses
YsKQH6ocPvkhJfY9SqRN9MGAUJw0tdjmwBtrsbsBIxmfEGtwjzrjp9a7mYm1m7tU
ci+kw94tFUKgx3mCCND/wyVWvyWCmh4oQR6npGSOhgmwQnAw+GwboGMElk+YMblJ
/k78lbTCgv6CfxeM8+BgAQvXgM6w8/gOUTZL7RGb9aPN8NlQVmZVOOCXip/utE3W
BNbexehy63m048xVXTWCRz3bxo8P9SxhcG9UsI2DE8/1fBYSEiqM0ggxra/cnib3
EZYC1t/jMVAj7284N6F7XUp4nOzUCbouHkzumDIcyyszR3dkeaSKfHzwuWAgcLHc
27D02ffSsdfUW3Ze2Xt9SPXTxcOGG1yIIgcgEyd1XviGscOMpy2drBOVN+QScVeJ
R1/xEnVdYPSF8wKlG6WlRTeRBtJosQvqDmSTTcnbnnaSsqM8Pwc81kP05KQKhyM2
OgyFTroL9Wm4dtpSwgoPfW4zjfU/jkemvs1G1D/CGUet0G71bAukGWGA8sMynLyN
A8GkJRoznzVHEs8mLMaI7gXm8rJDmFAih03QlLpAHd5IG27HdCAcF1k6eRxmB5Gl
5+wDqvNu/+Qaq9UBOAxJd1xaFn0JSpb/yABrGB397jnXxvT4Yjv7ZDOApCYQRZbL
uMtm8cSHiS32EAE9beB6JzWdpNDL9kkCsdKoPYN5+jwrY8KYx//u+fZ7BVYQNhZx
C9/gL59fJHTx8yGiPU5W0kIpWGjq68NcRWglcfZsBSaFWiaYPkn3xRgFK2Zp3cPe
TGOTBtYwkDd6DmzT7SCdQ/yAYhy2Q2mJSwtSg6+VQHgn4l/xVW1BYqxzXpZ+1GIt
kUzX5CRsg32erHO2x1qnuyw8qhJj63Vob3h37ECKSm7GAu33qqCfO4BRboSQWBja
UwscKdY11FOUWzlcnW4+15JKXh3X4QThn7buwPw03oZOu6p9XHXRfuZaDfEIG+1U
T4BqfUdqdjD1Xk+q6L5JXBicKV39PwDeYCGyy1Y+GwVypVWFCBi8LxtMqlUg849u
oCHP1SRSglg34LYC3z3ScDfSvcwBEx6OnLzy3UGQP+3J7PWKlaWWeOP76uHKolEX
a088wOawKJ5WKLKvE38Ha/k+qR2J854AYkl66U0fUTYl1iHaXuZ+ccGmIi+dK9hC
eDGxflqe+DyVXcZLKmL2l/Dop5qRbWA18art7RDWRdfWWbEJo9711KewamxTaeGV
TjIgW/9bbIjYsHTqVjO4s2tpbtdsNdH5ZY7LKKOmU7C5Y7ZacNdSY6fx3YETDZoz
0J4AyA+iFcK1LcurGCIAldUWMuuwoMFu3Pfw1QT1LAJbuzv8mtUUw26jt+sQOv1C
Whq4c4VkSNIAITn1EjW1t4NTXYEzOBVYFKLAWkgHRKVjyaeUyxU7x/7eR3MEmQRz
VrDqcyOjDvacjJ9GFHs0BK+8Oz1DONf9ZA/w5KhEWdLYzhTBL62BPw6JXiX13wEP
9ZUutLPzDTJY42s6frEUIwUgsFwIBgAEsIHUHB82c+Q4rksRHrVqRSMRhu7jGrT+
2oL1L3+zjQmZ5VdeYsPlFxgbvL+uV/sC1bI3aN65UrFlRKru869lrxzptU5i6DwP
NfMdpO/1+Ea8h+w6XNfBIOB7K2RYoDctGtbrWf9o9Bhj6vnklSKIBYTONXroo22k
K10+qyo/y6modSQo/t35cBJxpCi8isUzNiKxMH9ukxH3yBzXvltoWQKPRSTHL/7f
+pypzXdH24CR2PahOQgq05U4/e2oTVk0nUy90DfW4wx7Qn/y0zvnlo02Tz5YsSMM
XRbhRZ/lDp56HGQuZ8B+qAg7bcKit4XHlGM9NEa2SXvCHOEhfQ5CNG5BmxNDoeX0
8/yHPnqwSxEO46Sg2hgAoKk1yhJoreVtjfnpuG73tL4JibiOdtE5a7TRgmNUgqsn
KWatTSiYPyyZPCZolMx5acDX479eDR2G4HeAVl/kov8mc0lkU3k9jlC5TZXxIzyq
AOPYNxbCPiPyrOMbWtvoy+Xcr8zB7b1V0DrbVlRruZp9RylIMqdTn3iA5FTQej6d
wYonyIqItpHxHo49eC5LuuPaSWgzZEzPlgrDTklqlzJmDqLbUZsRRuLWY+isA8Sd
Loc9cW/ybf3frZvqNHTfgC9hG/8D9P+wdIoejIw8mnFICkQ/z6TA5X7cDKzQzyCn
ChS4EGmhwkVZ5kXzuiTBB4EKuPilR4iKT0rgCR/X9x+ZGJ4PaojpRbGTbM/DxMLW
wlTMhYgNMTnQPjTt4EAPzDNSVpQYv6tJzQHhwT4EqxElmLAdV+8L7hxLD8KIaWyS
/RsAwYFNrp+s0kJqyPZSWa9J17BDxXGBagCeQagyM1cBQKci99grcO77ukAEfzYN
ciE8/rBBDJVCrpX4xwl/6tPMA4Z+jdOSmVrFyTCIMLmClLbxVpLDRlqv/3rP4fWz
2GaPkg5lcF3h1bDcsbmTgLcp7SFLuSkZwVqvVWHZlJzqR+OAr6BQnWs6fS3nx1G5
eRDWg6w09hRdeFW44VlwlbaotYp7zFBfiAHigfLsZTiWfFQYD+jWwGdK7o98qHOR
rKVQlIiZHlMXTZs9618N2pSoPvYoCesDchcc2qoaeXSIOGeXPwJA7Oia9YyYy/zO
PKujO1r3K2u5TF1/hIkSGT44QQrqn4886zw/fhkrIgdQ1In//qCCfGdfDMfE0cV4
hR0ObME8OdbVqRsA48QLuBHojR32Vevq4SCfU/Faz9+TcNS3Rfg9RX3xUJ/ST8/S
58KpF2Yg2v6dB8+GllZFNIOJG65Gk3KPZtfxdZKBt16ChmFphl/yVav7N+u+huWD
OKq9hK6VwK6k5ERXYhBtzXojHn3/B+YwjkG75lIDDJSlRyxwVkFn6/lxseQeAVAx
Vio33dbNnrIpJ4B9UFb4mscUB4lRek918kCn5inCpFaRQ/ZMUrUWE/5WBhFV/RBM
1f13Ajny7iBgDGucXE2x1HT4Q7ITbpbFeWvDKIAFRyT8y95nHa042/F8LvfdanSK
pdNbZhGeb4J4d6InoO0dNJzlfjxRDrM1RhROgWbrV8TrFgipsgRPVrr2aKfXQPSe
R623bfRFZMyqm5QEYz+KN09PGkCxgG3FPvslB4qUoFGG96032MNYfMkeVn0hCNPr
2zUGkuEuzT4LJV6Ui3QyLTgJiL5k+fdqwq5FjGilxgraaVEP4oBP/deDysVxS5oS
Uc1223yiaRitiamLDQT1ydXlX3p6FuabDOetfR6lwrbMVa1tsU5USlloq+QXCwy4
d7i4pNIzSLVTppjA+CXe/TIZsj3pBCr5d8tg52RPyx8kkxsiUW3u6jbN2nhD22V9
dRIpR20EhBdL0CRq0rVzqqTGGLh+1BTBN8bskgHyFDa4V5M3iqgRKOifZd6CnmW/
Ev8QeOT2FLzkh2b5u+AzMFHXzr0t2usv/AI7SmQjYDK6y55ejSLOmxcKf2WqrA8W
sCw4tOgPiWTLZbfysxomr8cF9a2GxFxfLBT0uchA8nziDJqSmvqQD8Z0sB4SYEcV
y4zy/XP2+8zquMJy433PwuyY2dOUrymERTBIqD+mebIzBDQr6JKkhOTn7KxH27kU
wvSJJZTaGLqV8Q+Ik+SR/+X9teC5g7ssFfkLICVGZXBGBVFwAKtsZlzqvoa069Ul
GiardvFjuZRpz/naVbdLh06B+LpqvnRoE+hyH6sS9elz7MEWNMZjTQf6ZpjpCo9i
3JWAJwYbepKwPuMt/11Ze6LbVgKFszQ8SENiKWv151/hf0dNb225jsnaIiOd85jU
ZG9AYyf3BhlKZmlRN3Roe4Yr+aBkzfMx7/ObkOU4Cb1vbpny6Qhj1SZ5gJ/ySSKJ
YKn/O4pjwsoOd3Rz6ejtB7l6vnrbteD3TUs7azBnZWGdZmlVCnIc1XEkUwwzmYZV
eVr+uecg7jMlMjvmNtxadYcyz8Mal68pSp4U02ZJTnVJ/ZaJ/ZwjMVNhLtgNTKFf
p2E84vgkM5Ta3u4bABYAfiFJW5/mSVovcdA+4lrYeWi/eqrBmssOdsJPknjkQmAT
W9q5hiMOyA7cjPAlN/Y8lAndpDrD2J0OsSCbLAy1Vrvx9isIaZENMEiqg4hyyuva
Pzn0tQYqFqhjEN00if7LYI/ec/BYwmfttOrFpXo5n/vRgZHiT8ETJiLMuvlGmMCf
SYmXnUKvJYIsqSlN3cG3UsmdiLZI5z/xYIFMu3htzBqxG5zkNQNtTm6KEk61FeC+
XjlntX7Dv2uwABksrmd+TYi/V6z8ss4wy24qE7dMfwC1VfOvgxUmMPfaxtvGfYp0
W/J0fpUTdNxGVRTvmO5HIK1n7kX9MELSlEpfNeyKYqBYMaoMe4HpbiFYF4ERgriQ
FnKalCsX9R3RnOqinDptj39UK+ubkm2eYxny1EIewG6QJxWigfpokdXJeTzUQLhZ
VoecMSdlp6YlXWv+Nxzyw6gNXvvc7AjoD3giPJTGljQwEzKRWBU6OYr1u91qcHxP
+BN2D4e+6n9US8DLoa5y8bdaiO/nwMeRZc0GfMtwRYK8FqcSxlMPnoD2hGxqtNmV
mQ02nmhS7FBas4nRq/NIbSU6ntBxQ1/Zv66qnc+tk48zkiKXBM2kvNsfI5MNtlnT
7CBS1RpbFEhYmMTUdd5FuV/Q+afwFKYMmZEs3onatIWu4J/GlhuTSpNuh2Z01zUU
ZNY+ayyopsfAfORpsNagyWStfp2TbMUfjNRVEE4UZdLWDkaMcaP+uQCf3mlFBZY7
2KiGdRvKcKV9nXHfQcwSOIUU2K2lsYmrIwo99b410YJEaQXkJVGKanIAZpB0fqsA
ZBZ3AQ6QX7XYhqP9JQtbZK9no5tjwNiaxT3P2x3EYeYR8rHetu7y2whXeLRopgPJ
YjbhS1oOtwxU5kZmJIYZdK4G2SCyM+X+IbmI80YP8gJ+C95qEdlw0uIZKLi3MYrI
TYxudUe/0NfK6FDO4YugD2UAM+gDi/Ol0Jw3twNaZO1Ynyn9wyP8SIWNEoRMcYBj
33GxlGNtx9UUJax4awqvc6imGwGcV6rwjw79O2mVVwRo6pqDhxjIRpwt8do5vy6h
+7573huPFZEtYYmMnHV4i38DXv2EkUEa05FAGHzVJmsgwJ8DsXEHxxL7+0YEhTNJ
tXpQSFwZYHFGSvtEXZcRg6t/f6zOIEMw709g05fbOP8mQRcDMj9ubgBPdKh9KAvg
5/i1D4NCDNxoHsVIaKMLowetP53ecsXKgzUHQDCHZyLXNnW0I4YwrWFbZXi/I1L8
TThpxpBZksnFoLGkQc2HjtRsO5+EaucVx52TJNbUTIkVin8bh+Ggeujxuv3xiwog
6ayPGIHxvriZvnJ4rmXlDv8aBduT21R3+/09hiyKVJVyKntifeVgROObIQQDZEWp
MDLoWouaip0nfSir+lKcnLuMl1VPMQ71nbmBgpz7lZTA0ZCZeoOlRpLLmTIu6F/9
69o0Mf4Geewpcclmh4Cj7sguWLeQUn4lYU5C6cd6wWGamfH/OJSEKtb55/U+fzTB
sL/jtwP8YNy/6xBpSozzyfur012bJgbSncOxo13ziFvTJsBh+K6Ya85oHOY+UalJ
9ILojn+wYfKAu8dX4fcK+Qx+KsS+ypZ9IhCDP3CRLmT3lTQvf92ckiaKy+Oad3aT
Y7c7nUDA5eKC+Z4js8ofsIc6hvUxkFGnomvaYGvcwSyfKfkWSS/g1+tFFqbCJUpU
Qpa2DQXVj1hkwarVpQkTOCGPngp1LhTf94nlrgW8Sq5rl/tSmYfJOY5wWySk3m2W
m74Ag9+dbddz78kGX61bB0s3bOcdk5PJ1bhnnNX8IsGJZzWkJmE3CtRTuccVLMU4
sRZh8mr9r7YL1PNxZe0NckS1EB8bcGe0qdL4YfxddR14fs103gfnuLPsh/DGnlMM
5krcj4zBuIvZ7f0mevE7fYn6sMkkAPrkU1kIUxVffOf+iKr5xdmwm55LAsP/8XGq
/FeKk3su9gHSitwfty6zQXRHwnLBOMzzujlmwB9GXZCMHbmrwsPs6Cq6hgKe4LOD
3W/uNg2BK/c/QVmAITKB4WRfYKwQqXTfSefD1MUH/HNQ0wkt6DCpoE+Z3XGiSoU5
xFT4MsCHdpPkAD9yBlhVagt4vPChX5sSVwtc2R8whaU0PHfZLnFriqQXqJsm3HDW
ZEYdIy3OGACKAOQQxsms/b0HRQ6Rmw1OP6g6Hyw63LQRcZ4FkEgZhbldVSq4Wmbl
exT7lEXWAzAFGICIOToR8t1dtnxg/h+WHH+mBuVp2qFUtsmciVCtr/8QekO0i4it
IKyhgdS/0EiYNJmdojHi+9xirykRjFRTQv3LQw+HbjkEO+FSqRGZWa8TAYDwkzXA
t5poVfCDPyfmZQtAQUQ1yywSm6UyWX1ZLH6rPZGldTjEPZDrJHo6iafuZphxS3Rh
T2IqjjPl+rzEgPxdCaBGX8kt6DwgW6og422hemh1cVgPBhyDiRslgpz5qZ64TuQR
6aUNix71yFqNb3ee5TNtHSpRuG7feCXR+i0EjbwV9uqZrsd6Jml9yKMkBG5CdPRd
KEcxaSz05gGJa1pbJCIByaQ17qQ51ajirGQ3lY2s1inEPt/DKi6u6aRk3J54nxYC
uvgGOhToi5XAHaDxpN/pv0e4SaDYkmF6C6LKRke3NFV9NHfEGoidH31AsxuRd5yS
WTUkNRklL1h4xrGS2FXE+LQvAnhkIYrHwj7r0rWZFe1rk3Nzi8abfRJsxPVmt2VW
CKtDmEjwmqpkrFzJT5ieqlG3xVnu9A/+NW9wlYc1Js8xCyxf2ZF0KYK/Y6OOV4tN
1X7Uucgw+VJC3alvdpK1AIb4eVyqYApfAyDWEfhQOmgr8QviUrMXRImwWn95pmYx
YnUTe71WP07z1dOSMG1Tjy89aIp5vLECmk04vt1rGnYH70Q8q7GgC4GW88MF3+LN
NODzNB/hDiHcls1UDDKXT2AE7yxEj7zUnNyioqj8rFzfkcFwVQ1yygbx/kGnQ2MG
1qpStAHuufeVm1xY1iTNYMvbi84ABm38ImRACWh7lD3cbj3ln9MDhhIW0hKSEtMJ
ZoEfjWEJd6y0Gg2xYtdsVaLOU5lK0e1zPSBlTEs5nx3deKx/s8QPzGLWaiDRYSNG
fr67tDOjolcUbxW9TdFXF2OhfWVdBsDCbBNVe38hI46FMyJyEtGWpwJwoG02Kxi9
UygkO4WpbC/qfNVcMm22hBfB5CQeAPWyKilZQO/GY1RKsVIrwU+PzsNmPQm5nSgm
fSOXMg04CYRfRupxaeZuHlvsI+h8fAzF4en2eNcdPRRQDCHBCHCCT0EETV0toVmt
7LPhsGHMGvtiGhKWYPF8bWVgJyJL4l+DucFZX3xhv6x/1un894nxWIbimdcaBIF1
CguDr8oQTiOqKjKp+cd3XJFDDpRvFQXAWWo0uf6jKf3Mqdy0pMblCTUC4APVpyYY
rADyTZPDMz0UdAsSJDwloedBvRmR6PKYiwK9v70c4IntIZ6uNj3rfkqJNcR7w6Wp
g/Juh7IxYs3uR5BeTSDHhXY4pyWsehIlA9NKmjRibRvboArB+XhWQtPhTBnO8jRe
+H9/6m5L9oTt7oTqyXyk6K4ACYlF7E2h2qdiJQ6O4KNoN1IMAZAxjQ9I00V9qIF4
a+mBK1PNkD0CPRxZ7EqXx3Tl2/WaVusaOc3biKa9AwaIvna3il+NAD5Fdnq5711x
ZaOR/EG1zqFclRlXGxXzCtkUkarC68I9TopQ0U3H5/AT+w/K0SU40KvvUQnPhEW+
LADMEJE7zFGiR9OL416y8tMW0azSkJILwO+QBaQPbXMzmq/5qIT+hKC1eP1ZpDAy
Vq6kd5PMaRteWZuPjU7v5P4PVKVzLwp2f/RauqeLs2c4JZgaXASU7aADso7uD0nC
CNak3ucboBRL1RkKRPDvFbgi/UUt8nVtsPSaCZ1cIWtd5lYAxXHaxnGz8+fhf68+
pHfkO7YjZJdDaRA9pkORTVAO1GscOh6qtGrBEHJTiqZUPJdM2R7bW/jt9w3A7I+/
R+E3fKTaEdP+sfyhe1ytJLUjIAzMlmrBOdZJ/PPHxBLWqlAOtn8rIygCLqiv2LL2
JimXhOoCYrliXxaBxsCW1x7bv2c3FPAu9QGf6EmFxuDclaQKPhIAKv+wHwEDZs/q
qQGxAMJaaXDTpyRbzhKb9tpOSES9QpyJFQX9iTxdgZ3HYZEXy5pXBd4qqaCZQJyr
pMmq6wbkrL7PsQ3QKV0F/t04E6674jWHaqMP/5PzfFWdoiv2jBUjPyf/1pr8HkjD
+KJ3yTcfAmBVOqozFmAJUCuD3qvmCxm0961LDFr6PcAp0CGZrs1cVnnJUbRMCj0u
pNQiWHRaLWcsowgoCqOV5sMgLT/YSkAzAha6kX4TABmA66ueiEZEbYeXu15+GxWU
hKvthdOg4KFze6VazR+EzMK3y/6ojgKMUzaBVgxDkNvoamzq4oeYvA/wOicINIvj
7ocSintj0bL7kuPGJllFs8BKISEJRDkMeIyhNqwPxKfm6F5O+1+1xWLnW0gpL5Ge
bGUsOlcbRaH6TeShUSf059QeTTaVVs/L6fMH4j1TaFJAbjQ6DNfXcRfgIp82JLCM
VJi/9w4T+T2tWtCXqX1aZsDUes23Dm36grK7dHiIIBSOCXotpY3LIb0wimkC0VHd
VnwMmzcuxVQn5gEnkFP4qDoVg5qzTB4j0qBMs6KpLtrDF5QKGxpHYT58OPyl7fDx
+QFHkgFliLSk7jBAUyWQ9Pm01cKOiPwgnNDh3hSjBIUcPjfKE0TuO5bIUHGlGyki
mDUOFior9A0Go3yyq4K4XdWfpkl4VtOfqLNY3NFss9+sMveePS3aYTy2ZNHIzbxq
BS81z0MGAKNP9ztBv5tc0tH6OF9Hn/59ZhOWsbYcq9aw3l9IAQmeL+dE7NwRkMx1
1Du6UQx4cNNk/radN1wNNJKdlZ53KZ8pMGCMYams15lCSyW8AAwn1yBB8QCvZkRu
PA5OXMNQPu1zheXaJwOGEswI3vu3IBnOB+RjWo1DwRMEXI+FOHJ0dTze9yWmQRk0
1oe7xS90eqtsfC/Mpr+yAcgioQvHQc6D3CcGbyq880vzwG+AnFQzzKMXcG3HUReJ
bPcgSvikzoYf9Zi98C0IK+lE2qv7nxwEml/1I/cfwtbDh8uIbCn7uvqx2LG9Sz8v
ng65K5aBNybEnxKM0JNvhKnjvBXSdNgkLmuggAVBFnloUeZXTOCRLbQBZnndHd/1
pi/c7owHNRPD4N0i3c8GmAVDdHQBliXu0iqYMDHs5GRdsZLcQ1LpLT6hWkQDq93U
62SCfdDbuSUHTQRDZrv6QKAFEvnNaVlwPBRWv0Nd4Tmd7a8RwLyLjXfniWhoeim7
0uLqXzUhTkVdvcnTtfvg58xSOOL8wC7vAbD3iFSZgucrUR++wwQDgwBbr6Q+1bSJ
pstGBMgoZyvAFtOIt0sB41R3Ro56kNtNrCAfrP/sPqHfk3BCDDc4pcwN1Ade1/os
GUdvmwJa9cldtLqGjs8AEHAYZrIKfwbeZXiDo0Hu6XHllMWsPD3tEsn5IawHiI8E
7xacq8Ez8Fhv33i7N6CndTPhRewARZw5LWDRuHaRZQOwiXKezZZUEysOlNF1S8b/
akOhdHzwre/swSpiMCuDIc/tfdKElzOwrRt6i2/zWF8x0jF83syN8EELKCi84Ar5
6Z4R56FRU31aBCGyNZOqke/mNC4tsrdECeg+eAslL3HQu5gAwsnTCZ8Rcaj+OaLU
wY7DK5ezTjoFgsFBsEragCvNHZ6M7xE2foS+k7PphgwuxZNGviFRWq2O6EL/wQQL
6DgSk+jvrMZGkNwgqFllkjbch8YWngESpJdqqAwoy1X8obTp2msckWRxbNLsrNWr
bwyXxLLn+3NW+0KaghChdbLMCgMAMmrxMLdlH2cuheynM0O5eFojEyjAiiAVyVQ5
B2vinbeq4SiVgivZht/DG7z2F5iUozWJ2+Yeiq65omixxADDbZ3vKBLaosgNEUyL
6wtJcyDC/RD0UjsAzSrtSppnq9T/GN4x0jIS4cnCrK+lGc0DZQVM45gVxqNFNmOV
a7dvbtXp4sIYxnryWHpsXYMcHiNJOcnN+n23TtPohJTKW9Ktu6hWCgFOpL4ckyK9
DtmeRYRmLhqtTCE4nzQbOsDZZ0LZecXOMxPibEWVWDwNNhJ5okZcBngivZbvMp2Y
yuziMxrnGCp3ibiDnbfbwaGn3wgCyMqmjMc7LeH0PtbFT8VpXE0KAWnU7VRT0feu
TaAtXuxqPbP5/O83aO052yMQck0NR1+wTssZgOfYi//qzQ+KVUeza4iYmt9udmsT
icbW8eH8yl7MaEwVaG6xvOJpPfA9ONhroiRaYSBIg2tfV9zMnXYOK7XPExX1euIz
gZdl3v0VSSmYkMZJdHfXSsJI+y4cXaK4Fimp0l1C0A2rTeEqVISgqn2MZe1WOR7T
SvvhqiWhgm6x93IUTTYof5+WonEQXRbwLOYyjSDsezy/CGVbYOVSee2qegT5Tjtm
ne6r50rF5W8kENRk8ehUPwpzTj+NShOjbeq8bn4SC9pU+m/FLP+Gl2TbxjoGhpS3
/Mpus2Ew/XiR7yq2g24eWA+1P3HUHY0gcvmgTPvFT4ik2o+weOuj6GWlPwJjkYOX
XAFSxxKor5hLUnp/W+hEC1/Ch/i8SzpkSu/L3C/rY6K1BGS44hbE8Coou1uSTYHE
hogJkZ+84uNtlsWfSq75QdHe1oNQjp2CHQWEDihT34R85hsjElLwMyRfz5NG/XZi
pndNMavcu0frm6vmuwtA9AkNguBNvpFAq6PqG3No3hTpQdoPTXBYBWBU1nyrHBgz
L+R+mQVDTOR/2z7RX56AqnfOdbAH9F6CVhVjJ2V37yfHlhN9hkGhoM5QJOglpv4r
rmScTg5q3FR0VAbbom8rYkJfFeKpzeDpN3zd3uPXwrYskG9QMjEspNwAPcP+b+jO
OhKSQChs8VNTslmyxyJDD7Ieugkr8JZ7eId8uAWp+uaAV/dGCbzIy0taSSXwxARL
cFSa0q17RODBTRzdrV4KRhZhJomMYKR0ujcoGVClIRG/X21rSywaiVWOgtJGZLN/
TqD0+aXRCcliHz0m53GMTGFZWtPsJBRMtVQJoJRln1Ur+nk0iZvTNCj+P8DrmJuy
wWZbYB60AA3dQOa3GagHYRhMcp2KtYfScXBmdVWo5dXEdF001qPRz6/9y/CCqDKH
PdLcDSl28OiCLymjVKUOH58oZlsVtWznxxUQnqXLtmDKOhnXvymeIIeEXjtrlVhH
Ie/YJkgirtBWXuQJB4ULfn37yR6HjY2Wr99T7kcCq3iNeVzI5onCJRy8vD87zRAF
0UaMwSsWbMHqA7p1xVjKNliKMALBwFXQ2QTu8eoMs0U3vNvFhZ+NLFSwBnmSYFNQ
JCEoKTbCVFcG2KC3x2s/psd9vpIpDU+C+1NX3imV7aIHhXCR68XW7PHZsfLAxbBK
mKOzTnwHS0KeoIGZZiUGNw18GHYCD5TlUmgfQtEbHDkTSbtADPItOBM/p3S0Tip4
5rIPFjvwffXMar7J2m9lYuZ6KzVJkWulK3qTAAsNWaO3F8YOIyeZSEk3jXiK1dF3
585dHRDYGZYjJ1bI+xl6LdM4V/doApwuu4FsK1Br4EeGrgYp6LMTB4UxbxMwaLcH
08KgTr5pDfN21Jv4upje1SfF64WpBHGPveUS/Om7L+L6286zS/guG6NEFj3WjBkL
sna7SbBSiDidjXigiggkFmlfPlhZcrh7n9wXx5rJpptodltnH3BRIRHY5h+Gs/4K
60kEIY6cw+pMI5nZvbSRV8SwQzJQqAjHy7DZ3R6H8x1IvAgUdKd0VW02vjskr5ZV
XQj3NHvFixVnr1wYM4uBJ/coZ8wmMPTuTPVDx5bFGLuAB56reEn+l4haqEMYdFa5
mWUuc4KYlOSePi5+h30l85HhlzEcKUt0qXmDXEIr5uIDF3vRRCk94mf3qRQMR1i7
p7fW35d1RaTpxwEaUdH0nOoX0SgNC7D3sYa93+AWTdVHAmeb23XuKyv5rRd7CAX5
jIcd0s2HPzDP6IvIe4sZbKH3gmZLyVA2K+tOyvd+Ky0CNvJkccMLboZcMM9bfxfo
rU3Q+M+v2kiwV1IITkn7Ol8tcVbxYDgMZXAd8/8TeIX3xL5Wei2YjQ1VSMt02sll
hYWiD8ZbU3SCoooKI4cZBWemtiyJ6MUWMXoyrMy2elhHmVBsXgCsVGBOr0GLiQre
dGTvogOQMyLg5uA2y3WW5UC7TF87O8Kln3zJfs16/4d7gUcnBhEJG2QuSG+fT9Cs
7H2hJ2k8ccbi6IJMeKD6jyFthhUpQ9cbUhrGDmbKgqaCbR3LDT9jAy7B3/7CDyWJ
pqmqLYgv2R/wljLdwoFzp4sS7fu8Bj0MoaQ+sAlUXeBxg+poT3a7CqZn331bu6rV
x9GrghT3JqWJrFRarcOISCHAShGPdT7FVuNmH/UCzyCl0WmDmXDMoFSk9o30LwJS
bANoOipfUMNPiju4qVnwzEiu6jC7AJgA53RpKkzaR/9rnPIVmiUMeTLTYol7ec20
H4Z2g+7hNUiJKXc7YZGvP3eUKr620stxdbmzZN4iWrf2IX1u23sGrbpuDLfJ9qPF
5AI0fcttKz8pNqHCETpj738r3CqlZ+SJk0nGW4V2izcn21jEohVOnyHtorer/1jV
WLNtOhbK4tD2VbLAbUfKNmenieaS13qRBQZz96pkO5oBYVr2glhW8IntMQkWKpcr
IX8rgxIBO3sH/AfEjVxN+x5/Dlhb8HHnH4aul5uf+6Cjx4uE5OcpzNNsdKACgsc1
IkcdQaKAf+LHFqUHGZXVkgADnV4OGFDI9FuHQQ6wKD3agt6+o7kn5pjWvyDeYF3/
KIMwmN0pG4qQjQP8XVnnn93Gk07nQ5K3ME3pyd25UueU5b9CsWh1NoBK22s4esUX
dkiIOAB00FbmIxvcYM9R+Sb6R1UcBfYa1iGzoSa1p7DhKqb9l59VALXvOLJljm26
dX3zV3XM11nrTFCCPGKMQJ4wQierTAYLioAFd9AOYACcaSIN4ALNS/GL2tuEtd9j
BxZ0exwFmcivy3m4x/PYTNUuapfAxTPk5mlo0Th9zqozNgGuNP7zal9zwYofhgZ5
Ra26qUfQ7bqWBMIu1/ej4rD5KqaQOcqECLK2z+XiuzBqYekC5/pAHmbxMu0G2qOg
JSkFjGbgWbathJSZgJjRv78fmntdLXN3y8qpc3sAkFPs1pmIj3KgWiQpHaRkuqGj
sgnih3PLRaALW7ozFpkajc/Rfvt7zlwpG+tnxXgE72MMDm5wysKo+Upg5QALixC3
/JmjB1W+e26MWWNoEq/jFudqXsDRT80hPdYd+VrKiJq1r0BUqrG1SR4auIa1zg8Q
Hf8RghSgGUPqeUaH6L+hVddCGJ5bE2/IiwWL/0zmumivvYytGcSt5q9/DB6LfQSt
p+uMXMVouyAeg3jGQS85wPMY59imUZl79RWjlEGKlaGQbto+0S71uGgZPR5PNq0Z
V8kDY0J+0GYLc4/wAj1My8SsijtOh6IfDEHHgvdejHY41aDl/dweq0BRlp79dWj3
3lSp2gG5p7U7gPyrN86I05HqmZvh2RLcWfzxshGwzUJTG5JOV8CsIWQtIkQN58l0
vu0XkrESoRjgp1DQh5LbKAs5ur58iqkbiJs6NMmgWY6lT5UWvmZCFcNOxXykn1Nx
AJlE4Rv/bAFCw3FYeOLvAv3gR6Vf9pejBirtB8CvgclIjr3Dccz2xXJS90RP8cal
6OZ48sOYCaVSIAEGcaMQmrehMJhhSArO1fvzMFvIbuqVd0UXg84ctbmcw4SqokT5
IP+20VhqEAiT/+G557zDX88xBWzfqeBn9LbSlmKxKJkKb7aZ5F7B23kh9WvO7Ik0
4BuTW+XoOkbc+LcGf795VpAggYeIWosHhhWrHF07xrQ+GXeLv1b0G1mIEwsiw6MI
jaf9t5n46UNRAmV25lAxn8SUDGz4rnL2y5RDuqG0XN4bv05ujf06QFB1O1TB72qk
h+q7ZbE0n8Tl4qL7y4iYeiFY0xlWJzFgrJHY4MBQvGqCfNaEWHvvqsZCW7XPPums
S3nsuNj3DeZDL1MwpV1JENyq+nBNzM7cUtskC9i3TzwM7OTKlHNDIQFwab9slihI
BzX3oU52CTxEnWS/aKthf/RtXys73z/svpNfwjvCzC1i5gKV1xxtQqKrgZiYimGB
8rKMCR6pIFbM8tbvnS+oW6YXK1uj8mVteWcrAejj1MrZNgftp8mYpJX/8Bk8YOXI
pM+VHYlkNKEkapfbHOyq2gLl9iNTaacbjtwPvIY7xZNzqWJe4nxjxxkzKNJvHZY5
jUvdm2X74aTa31gI93WkLkEheclEo/JHnF1cpNZA5wggBEhsCxsRhBIPlHLCHd0X
of0nYORVPuS7EPcw6TAz3hExP7FE/3D1mJ20FlRM9yOwywKIRbxB5X9MUBovC/fl
9MxsWAS2k+Ay/unCfsXs9T8CqtIam+mLx/rs+Tn8YI8B+7/Dqn8Py/eU9zy71489
63jbCRxQ96jFcg2tysiZ6yxG2+7u7AykQDafwcGRT7uEAknSDYttZgtlQrqa53bH
7W/Y7dFou/Cn7nMcAzV0M1u9+ZuvvvqKuJIBKtoMSmp7tzZ8PBiOnSDbhhzs+Xag
tzQeJGjUdShl3hCVJ103MnWY0rlwY0NxGGfbUahbrOUrS1nzzl4tue1aGJFMXpG4
WXH11VaREzOKZmBDcqREvwJpPQ4DLxwkKH5cPePySF1faV3U1Gb9SW6w/royVTYE
LNCY0sJ9un21vw+KEms47YrthAsE5N6pmHuVz8HlfUgk16M3CP2JwMGToN8vpq5M
lYZaCSO52HfTbVcgh1LKK479x5BANX35RCGPhn3uTARWswza6LMT/k1iAHtoTkv0
2JwT3CfBu4o+N9rIxj0LwAvczFVPhAn8PTeiG8Z77um0r+HNbOtrwteDV+XkRO2W
NLkKq/Xw84S+MfOGXDo/lqtYYllSYOxu7H7Wo6KQdtcBq/rbjoWDEBodQE25etlA
CwzWm84ujnFdMC9r/xkaQF01NNFbzQnwXchaGKaoWD4jTyyl7KVp3fUpxDZE+gPz
bzAKtwJQAvCm+e65O5C3us7xBOGbu4lWJKhZUlBnOjmTfizf8bNkvrsCgrGQZ0e5
GsSUbGW2KenohFt3VVqe7E0pwu3c2VXVuYONWfOnSeK0unbm310tgkGd4hgN2XqS
pPcg3KAMZcSOQFLzhFfEIdEsprHuZtnB35YhQvO7ipjskdr8t4PEmsdy490HxHms
pxlHAh5qSQPmvNEy/hkCXKkLyK27pBkbxpHVUfUBeDWLrPR62D18jOP0Pxoeernb
NZoV9obpt7ysfenNLzJlYmx7n1l0USz1iLSe0izEjLO/+YrstADCUZYMLwcLySt3
+AQqfJVlKIBF6b4wdpwH3n7cjwyRUOUqLgNTd0EyCxhcsDqNpOV99gx3TNcEwB9H
/drK6NnHFpU4Jq6tsMz/6TYmT27jR37CYCX+BHsoAxcI15wzhjfsET7MFVfs6AXW
tVbC2chKlUduOGfPnsfkoVzgK9XjiLt8LPdDju30g+syftCSQy2WPkm8dRWxjHhV
vcNxgQZAUXgz34AGuGL3LlSHHh9f+LSojRfvwKuJdAccZKCL24QpNpZg2zajpzex
VRghx+P9UDdJwLsCXrFbBpJVQNXh+8p3xledJ9kac/iUf0buAp/vJPHcYXzsDRKg
ZHDiHezfzZ38hUgUUYZ2YjpMQSaRkG1WqV3yumK+qb+nM5lNsaY2tn6EAKD2FWSr
izTPr/SxTYRj+13CT84fDZUaxHvxHvv0juuZs/OohFNg05Sbr+z5rrlOYr83aOq6
oJEMKN4uRdE4RShqjFrimy1a4H8wNDHaxFCE9Uye5MgnNX3mimkbbc/rbgS0j6Ei
p0o6C4eptalN6gZQ1II2j/VI5N135i7muyU868SrK7RX+cCkGYdR611nqYBNchmN
8EbmUwjLg7Kt9p0q1YC07o+kBqxn6HV2BDkkMiI1YJmGSzpd0I6Sc2sJhQPlhSH3
owRo8Bb/2Pmm08KJ++0ONdlJtreoZHEUZ7mAYw/0WWiASZg0iZCpc7iGR2+ZDW8v
hv7gbwUL6C2tJiAblPub/CHTfYGG8cgq1Gu3eotPw+5ryYaF+sqaGjBfEP0cqOvH
9WrVNrRB+BaF2ka/UvkGYeFE5CjhQtqbmOEPxkI2h7I3dgbo/2ySPydeT5ys9PCs
GkxeFeTuQejhk5QxvPvnjmWwuTjwBGdE1KB5TJdoTJrzu47mDB2htIrTsXrpwrU6
ZzUYKcILldf0rIKboKJjMq4tImJSQ2XmWO9Cs2ioEtbkPeENFsVOAk6P7mM5Be6g
Yohd79KBt3pvbh9I6pQ4lWnuzPyQZvaSlADK+3CuMTJKwcjIZGxJ9tPhAtDG7c9h
hM42MOGOSTR3K6ANVPIcIBjCDRsnPBEjbAFEoOPebmlD7oyTHpKuQYNYHmCY4tUH
Z0mFkywzY+z8QxNrzQfMzRL1sgXxMuCmFxjpFYLJC2bUclqH3gj+xcblWkwNrBU7
UIPbGjy4izs7TSTWjNxFd4eR/bO45zCzR4yR63s2PodnOqDTr6MbZHbUt+js+ajS
9HFsb8xUwLI7xDKsMJPpxPqZ28+k6Qvt6zKnRi6qCiP49nD8STgklpwya4cF05oP
urmKapZ6IzIJwcYiGx8JS5HGBgkaC24rDARZDVIx62brXb9ViAi522qN9F/47mnw
BgIsy6vgw3ZR+ajzMgnZS4PPIIOEabAbFMsZH5+s1Kc7zD+ER5dcfwIXMzaX+jHj
9ZmlBmJGoaWGd1N9RzxhoYqGNESHO+v0fqRCcqJ0CwdDTeqRlFk8nbJ05WwR+yBt
naKsugNewKCVfmHHpTkg3dOAuu1Esv02Axa4uCk/YrKFQt+oxB8a7OksZXbCH36V
bokIUF6uljyDROgWhayalpR8mvmqSrj1Lu3poYfLA14rsZdCspgsRgDBasfsIqYQ
d94BnsJgRqJO00ZBcJpSvs6owVeYJjJ+aEC2v3rRYgapR07TqlREOKYjZOkslUa4
TvsgZVUfmvf3Wd3QOF5EHKMPmqLFjZaQxWLEgonhgA7tCr5lS73KePm3wJtRP6mj
ZulQi9jLBHjW7qachlNyIWLUQ6sHv/FnRFshKV58wmwJs2Its7FC+eWh1Lh7/Le9
mCpDnl0tmnyjiEIvJrgBWg6+/K/mq7F1zGfkTQTYwUJgQm+d7/N39UIE0D44Dv7u
eUk81QH5YETVoRwsHa6P3zTQpZFvVoYoU5faUUWtLxCUrwxAl3jztUPOxqDMKQ1E
aqFmlsPlw9DqK5WYSdmqQCJ6SSvZgbiGZ7+WkxGWRTC82aDGJq7i34EAHt/8jaXW
9/vI/UsJlP1VZVEV27P3rGNoPocWO/l3i23auwjieSm8VhosH81ySDHXYw5q8xy+
gA3B9lHjMeJI6igAATche5nE6jfjpLs8+iyaQH/kA4vUPAaR1kgaTPFlEMxO+aHe
t9VGrwAg9YhKm3mkHd4PwY8YuGhwP7W0vv6FzJyUlzbWgNsFPqWJIqb0+Pq2IRg9
0o6bFk3OQ4aDPSLIOXzGOiGmHtOwED6NRTOt/awTrSk/PeBWjKfnS1E6Dyjb3Mub
tuhNQPlfif4U6apg6WkcQs+Q6B72+OIZklivHrOElYaRSIA4GE6VM8llx3wIS02N
oOYFR7xm7E2flYiN2LIUgbfgHTij9VXCQ7KT8W0mIdPMgsIo5tKt3Cv0icUy7ga0
+Iz8fTIDc9Afr7rrt0AV1z1oQRXxP/1Pl3udkrT1f0P0veNQ75iX7HfRdKM9x1hk
dRUNwOxUPN2y7YgZAN8edWvkwsxu2zyShx2x4lCv2TW7jMsIQv9HtDqCzOjczgjf
iqLwa6E0O6XEhYK9wW1jPfT9jgSSvp2s/MH2cY46ml7H7xe06yiHb2Ce6QWECza0
9k9ozgXEJltKnkbhhcFBaM5jGopovwKCxum23lfC37H46Jt64kKu0fJOBr+pN4dm
SkQE8DE6HZsoT9+UeQ48vk5D/hXhbKSnDPSJIwL6XS5OUIP8hLhWWmZM7yf8F/7c
i9LJNxyzHJSjZ7nR4ixda6/hZcd9y/Ewk/xOd3h3cTaMU2/XVmOP1wWgwvhSuEr9
SXquBlfjpzGS1SS0dtgV7WIneRbQH/9/SbRlQnCp233cIOFlU1Z98nBW+iCZgkS9
G1suqGkdKvbV1vNr0hHXlRqeFLPlFeEBkJXi6EGvAo6OAGQHU9SaXtYWdIGnjHV5
rjfMAbfKG5e/o1Nv5eECBpnfk9ND2L+oSWULXiWFEUiQoPA47cQvt/tnzZ1+mpZb
tVOpoY6oCefDNSvxsMRjKDC6O33wqcwHBYCMHfFYs5WwjjirqkY0XKd6SdUMlWur
Jd6Jdxc41ZUAgf7x/qW21zxEcNavpZpH88jtPIBaj65ll9Zmio5fQ1mNquxcL0S9
CQoJwmO3cxztZahEr1vXCsC5YLvjOs9fqUEZNqi8E3prN2LCHJVOKNhfrpgRmax3
S5zV4AQUOJ1Ss/tTHiageqDwibzvmuPmbpm3qQ97TpzLEOF1QXHkxtQZeMVaJFHM
JcC3RvQYGWYsCOuv3y3D5Jd+vVQ8qIRFzjtCs46fheG76qggWAyQfkznfJ/+Hqv7
MFMl/SlfXgm4LH/EyRVkJ4MxG7cMey3wHz0IRxFi4HsHnv1NEtmaChS50dLpue2G
a7Q78Ut14zNZDMKQd3beUv9Bfeiyoys2q/nVF+qFxdCFmqxjld4u9UXaf7w/0Rbt
mXuZk4BGJj+sVzdPOOkg0+G7W9yg9lNmDF/pUuldujMddCrBg/XdFD3OT+AK025j
fEFFI/c9w5d305CMHOO/fEsBFDl9Ggn0jmU2tdRJa6VR2s67Z1KEnn0QvSyujDbv
leTHxuYkwLnsGZ6iPj+3ydFY8AOLJPvZG+K2Y4+ha64wK7g4P40P1OgHzhz+wh+l
QoTm5v/hHwN1lHlMrMarYuGMeAH/2FPOwHGSBO9Q0fR8R5l3rvKjwW0sW/Wvj4UY
XcgJwo0rNT6er7yyya0B194MuRYRfZkwaGOhdSdmOYENf2Mi7eXlNKtd5hrSBe76
MqQKrQZwOl8jkWQMrWLZ4GaO/9Kwrr687i4+MnRwYU/Yuk0zPkxan9U1AuOni9o/
FmIzW3RrUg5selHdMx27BZfI0vZVh8SHyNF7lT9vFaxLfrZFSVaj5NgAGA2tPhH6
rIvk5HOjVGsy2Rzqa7+3T/dk9MxTQ9VFUbbieIyMlZBDsoTcW424Wp7YsthK+aXW
lO/9hlqkfKxZl5GsGwfQ/d0yeIh4qQ1giN1A2xc3OmUSRCcDfgXq2YmEcZT/tAUp
x96jr3p2XYxK2yoEqX2LuWabET687usbGMP0JdqJjcRQV5zuAlg9LwF34ufpLNm7
Os4KUgDXVmG+a7lqML5vxCYx3nCVlSn9aVW/Od72jUz4aWj9B9aSw4+XIBTM0E4e
NgEQJntaSS5oqM+WFErckyIKuXoNYgK21H4Iz7vNfY5wkvQcNFx1o1/QviJWFopV
rprsiN2bcqvO6fWOze2qeYhhqUiqTcUmEn81IyOq8hWtaLXrY0UiyqJeDZpAQ9OR
PANCJh1wP/0R79dhGYEeSYyT3VdDHg9rAqhUYFlEVAuKoWtWqDKZwoKkoXkJNqBr
s8H1M05HHLvw5KbB35Gdbxy1zOtxtOJJxRzEGXfhea7gMLHIxXr+39YHqTr4Mu4Q
MVutdeQ3pANZxOA+mTvnVb43M2DKtF7NB02AZuGEMdYF0h7vsuXgd6OLUh0+mSAE
Y3I2lTd4cLzpjbWRI8IWjcL/E/BsTmwxeC6VnE32peu8cZ8AQTkSv8xxToh9H5R0
YsptL8VxkshJETq059/GJJywrpT7iMVja3MAFdjY13pxnCYfPbgg1bJXVwJE5Dud
RSrgsepirNsC/7wt9yYp3kz0xRQQzTFbT42S+ZB/87ruf7z+xXB3jvuuCWs5hAML
O0hxo+aBBitdnJLpQDdczVQo5Sq2EP51QwYXIDHvl1r7j8hGo/bSwWBb8rGkpkmY
SjiQj0BWX1+CSwmufJXh8spzjEj3fCnLIrxP9xLKuJ0Jk6Va6q3rkl0pWoiE36IR
JDmHz2UM+IUve86yWLBJUdrH+xPVndmlX+s0z/lUtxuZrIn9Cw6Ncw2GLN0CZcdb
52uQf29mdpCz2cdDpRykPf01OB39Hgq/jRoUHhK5SmNTgoxGl0ZrgBRYTqxivJfq
5ZdHKJKShVfAs4tBCccwfG07AowHUctPMXDtREpIpqtbRDG5YayKckQZ9PS5YZCs
MMS+gyLNDCBYXdwzfcoli12xy0eD0mkRoNFvmFo+tf6Yfqnpyb/XKb7M18qjXKYI
H31hxNjO4oIfjUTxxju3ZRz5Q2KLqh7Lj4Tbegm+f0q1TOEr22zK+NpX5ouBz/0h
Rk8XdgNHtj60O8T3lZMpVseR9oydyCq+oP+ZyCbGnd5xseWSOcXD2kxHbd341Zuf
YHlBvu19mkAIUhqCXiQDG1SHRfNVccARXL9M1RWCOIoBpes6UtEIlmn363Ipa7hb
NaH0rwCQEQphzV0VvQ0lAjuBslJ89Ir3I709O1P+ZbS1GgUtTueukut5kyQTcNAz
hJriHgLd46+MLycEAteIiFlCC5MnQL/nl406S+xDJrfEaZ2FGpUHl0xy5SlnKgyd
+OieQEwUXTHDbp3lMo+nReWicW7lc/x8LCWfuxoO/5NNoeWa4+tAngxnFoSQldhj
JN66WbjMA4WOa/ywkKEXD4IX+wfbkFtvkRg1zpayAhpIaDTFw60epWLkW8PsmUQg
EFFxFPPq4tsCRYjxhJi/ZMgOP/x9NQ023qUVwk+NpS3Sa5XfUPKEfsS4Le3WlZSS
zQ5o9QA3LwW99lgKBHr9ml/4t6zyKcYBhxxUQomLA7jzBIQgf7tgOHmwJl6/h0wl
jxqr1YNkAPfaP2jVasgMyfsUKchUiQqHFQkeO+WlVvqC6IjOWq+2k7qoqQtJBrmR
Cpt2bYYOlbTvUcy4az82lgahiwVXjG6mr6nBkrgYkQHzgghhMWAvDo1/yWYO6DFp
Fp/HWWMnov+0J+33METtVYN0g2PzYyQti3sQ24XZAPgd+pemgAZaeBrsxWOj4D0D
WVJ+AfzX9EWlVoZi9GmQLpakG3nPaKnVyiKrXQds0LzRWbjZXkHKqUkryd/Ishc+
HcSnDQ2t4PlqRwDazc94MY8zWQDri//+3KaUFfER3+KBN7JcnpwGEHfYEiyuQZsl
vP7dnj+/0FEmhBhVREJOE6EhNE1RUv4f2MJkoFUpn5s864bJWPlh1thuwnEyArLe
GCpIEw7yI99ejt5JkmHArspS47CDRPsj+xqEFEFT/hiR/TTRowA2zmmZzJuHAVj5
V82OUEzQjq0DnXOtE4tgUxZnYBtWeIZtjAOnitX13snKOhZu2iD8F4ZCbEK8XiQy
+8kHhRB1JdGWz7SkY2Kh+xGmg5OLwtzHrGgbYjE+QO8BbrEVIESrvF6a3d8noZTH
IizvBL/yzDNbYPJkPdk300HyhYrMLWfjVAqkTG9v9qL0smN10PxJaqfPl7Y62o9Q
eV7MyuMlv5Kc2wJtq+35LX5PMIgrtZKnqcDUHC2oNc2mhxRqD6kv6ocv3k9sYNVb
/j1UZbVZwtbfU6vAfJZObQDtFRHR+QW9Mh5X39ynZ99g42KvhQcijby2xneTmb3D
FHgLW2oA6WgWK7D+5Ek1KFQnpR3G8NjR2s7oM7vd9+YvVwSpCeCpS1xJhcHo99wh
fzDQhXmommSnmu7RI0BPqjoX9k/JNDtfaL1BHflOFiCNZUmhhbcAuNnu9fHkNbNR
YFF456hiu6QkBV1l0a4H0HN1Mt62M5ygRlOPxbHWCu40vS9WQkhl5bztFR/5i56T
auTSTZayDPu7jZYxpD9LmkwuD9pkAEFC/+OnkNscwd0BvpbDtpaKeSMz7hKdkcXO
wlpDgSSfQkbJeBQFVOED23BoJhJP5x0358UuJOWX+GLsDPbzR/oIZ78WVvPWjJRw
6Afoup1MbkonmDMaKTCQZs0NBKrDpm+CySLhGYTywaeAXGU1ZbRwAxR2OrOARm/c
Xemo6fd+VX7+gsqSoXgAgeIa7zrwRX7mFHy4eH8ZEfTeShyk01WadbB/s4tafoYK
Dbkc+qp54bFTU51wfEqDoAZ6r00R2povnRt3A9aH5jA+0zgkpnHiPVX9huRK75X4
MJP0q1z+ancQZpMbkAONWw/snFYn6CKIyu2+rdxlzJ/UNsJytcoGonE5GsZrQnU8
1ZmwBvXdXl2CSHPeEGR9oWujM/FhxSY3c7VP510095T5R2IPIS9phhc3Y6INjmth
/EmmbCoDtCarx86u2cHYTOevZhMV+04uSNWIMSw3baPmTDiZsMTI8jf3zz1m9+TA
DmEJ4y+Ntk+gKNRhgRRHRMoSk9dZfuP5I27uKN3Eu9fWB8Gge0+SDXxc+8GUc0O0
JYAhQDiaKrUi7BJGistEIuCXWNOdF7Kdg6R2977eDmpqs7WT7BsjZgIlvRb4tFqm
dLCCghHxhsiqR0pZtm++U5dWNyEAn2ONnkHe3H6VTvBonWbLGRSVnUP19ZnVbGlD
rZvOPpdDqQYe6GcNtUUCI8yqKY9kTWvkrfL6zkL/96fMl/whYPgk+IkVRDKL2Yqb
ejYc3rthqyAiEn10wGu0NzSdpGIOAe7y9ILgRSHtqjtgon7PJDoUQ+3c1ON5NyKY
h6LocrK0K2KenB+Cjwc8keSJyYfDEbMFDECzxaGT40rBSM93rcnuFHW0lN29pYhY
CTPQqgDTZaLXgP6zRcuH/j/eHFEzwh+s45FendkDVfndS53ZkehNx0wXh2ERSCuT
T59RFn+2xX6FDQAPXvaccypGlyyh1DyHSTPhH45n0CL+X9OjD6fYVCQNc/byqqTa
BoZBAW7eTTbbG0y7k49lvKXsEQL1PGkLcnF0vh1d/WOiYISZ6XcAWpEmi5mxarDh
0r4UD9pum63WvM3VjjqGMPVuOpZWaMx0Ehvaf9Tz2AEMQ3g+CX+MUuNcwEJ9e/AE
rYUTiexWzb6QXeCyYkgyoLCfL1J113xQP47urgnOBWg4QkU/GLrW7eRv5JQvd94g
1wW9jb5WwpN58Cp/QhZiJKKBwrkOQMKjoJwKursNMHvK45rph4v5rCKBKoC3M+ZL
DBUwOekWoWi6xtcFoP5y7YHrdDNIyeyonHfZAloLyMug4skEfTnlfwzqA1FUjO8f
fYWZ4mdbt9OoVeKMKPM/9nz3VPe90LAfYclm+h/jEO35dp2ukBFO196odJcfmIn7
96pi5KPKy8cXWOCS5Ni8xMSdVhGTKQY4oXC48qOiXhxqa9ruaUdqKprCqm4PUBAa
ogDOcpDtIAZxT20fYaOmK89xbNhITdlQG+f/rbKcy4HuRtfjy6xRUxf0tiZB1cKA
rPoWaJvD9hTWO7l4ShOMjyIM70aHUyQ/off/XPUMB+FukUggw5mAx7A0B6XefCRC
ebwCq5OsVIUeMQc1P6IahUB1CsraMAVU3m1a1L4gmu/ri7M27PzeTdDfnfdCyi5c
hzZ+8qtm5aW4B0c0MM+KJz0mV7VtLFXcTTbXTyNiWAjQoT+cxzyESqeX8ZuQpzfF
HgDbB73R0OMbq7jbrfIjrLhef6asciKGTRjgS7UP9q1TJmxhmDZhI/TERIzN6jMR
/CRp5HMTi4EXVl5x6KBxjyowgYyyrf/YSJmruk4+cVvD6izV3eWTJI4azHQuJMpK
v2c8R7r9snbygL5M/qNoZBuUPFEkkxJMSCU3J6OBjVQTsfCKmfibpVa+IgIml9Bm
9woiqoLaF17HlRsz1Y5QRf73+JlOYRJ5h4KlljiY2EwGtX+MceJFwmr2c4s1T422
fjtISl0Z+foQuit1+nHKd8at54tz1SeO746kLxfXlYAA8cE68wux7Zm4vSHQddDF
IAonW4tT8IyQBtw0MgfJzKWEGvvBQrPV/vpZekQjlWCkwKbNS4AVComyn5MRmfaz
lIOPe6CgEAh4XDHi4GGf9sZYqk7SDXT5VyvUGjrQQxzDKldnYn1gvZZADbpGKZAj
+t/HiRm6lpt3YVRU8b493gX5BzX7ayQvuNgtLvaH2I5tR7x3cVEKogEOSX1g9v9O
4QpGeWue32d6a0ZfRoJj0GSPeRDoB4vONktAqcDn2o2Ty9iAlvWxrmOB8jyEZZQv
1ha/pdOxIWzUPhukHPHRQLo5TbCo+ko1BHKMkWUYK7A6I3T8absKIbYw3IiAEcbq
ysRsSaoYy4GozqFIp3nrt0ANHpQ8sUVKNgUbt+YD7/V7ueeH+6IZTCg5649S5QFh
FV67TkNW6wGKuCvREFTRXp8+m5LN08VDFwAiG1itr5Sslo/+2d2/pZsw0kDyt07l
tPLnNuaCUk2d7fgquLwa1/curGwDZE1YhRHyvi986jh1WgVegEvAQF0T9ZM9x43w
xVjsmK4heq2zt0qJ/MRJ57eSC1Dkcm6NnljwQtUoCzMIV4EJNF0aQTCLyOuhqlId
86TuYk18gS3/OV5Sg/CjQ6bbmNH6r0uCLWr5hy3nmSiqFf5nG0mBv0ZT74mx+U5l
Mp4p4jZSP37k+yisbXrzmQ4d67/Nwqh1u1qMlCfyUFCZMTPfGEWAKgm+BM+3S1JC
dPNT22SYi40jdo2HtY5Bmmc+0sxTYEQd0XsYbDL/kC68CnTKqF5hukhXxGHp7GEt
uSPyYW/Ct6xTdAC8LnRAO1N9xUenC6X0X0t7jOOQ8+YBVhP8NUNL/CVV69HTBj4C
nX6TM3OnjLGcXyPAJyx0SUn8LH/Oe3iAGzJ3fixKPb3fZ/PFOp0tN4KrMteqny6U
0ZI/unTT44w41kigQjtoje4GShUUmmjs145Cz4dsWz7yPkGaIJPONb321qyxSo5x
9fc0cBsceEcKihh2vV0ljXk0tVbIprgeGdNcBLnTIZm+jgbhg8Edd6VrM1Vmj0+F
wYUc/ozsdqE0LGdYC6ZBKGd3mNa81pt2BFOCaZdYDq8XU4RYw2dsdCQaYBHx08nd
NgsxSXwCXIFl47BPFSCbbN5ju3LEJ7AStUFLwqf26945ucLXjLh4jTxVytdp1feO
e5+gfP3t2XCKMz/jrVX8cM1VBrbzhm069UiPpn8gHLkNVv688FI1ZpEg8N9R9at/
L+0NUHV18zrXaqR2lQPT9D29hNmRGumE3U4/eM31krf0vM/bVwq+wMYEkOtpLAr3
5aI2dpMlzq4xARJ1DkLe4nrq9BRPRwe499H8cjxkB7b3DW2KwzmwD5Prz2KfjX32
Vp5YEFebnw/mdAAoGRH9irsBbS7P1+xNkAu4E/33ii10D2DACiLXXtZYZEFxA/nb
7qUyWbp4dJOjUstukYZtLoz2Zxyzm2IL86aXIufhdQRvSwxZdLqMGxviq2RlUTkJ
G1DXO2m4wa2YhfC1B1Tl8Wz8Nm+8zbV4LhmVxaHaxIUNV5Di+fwLrSLwAcd0ESGi
GuBmOKHS18pd9jwefYuFwoLpSWDZcUn+Luq6rbDTmZFEyhJ6DMQF697Q3h2qsl9W
EtS4fBw/qbCcij7JsLmrAcNMkbxW3O7FLnnE/PgRxGySFvOnctDGYEM11nBCvxvT
R4k8pIVhb4s8rxv2+QxcFnVzz3VceBE0viIQqNVSglb0nYA+ONC9GO5IZSZ7EKgu
HQvcHyBeqR6g8IcmXcHnNUqtfuT7VWx3d43bdfXdm9zX013Fq65SR2uJoRq6UhkT
/jETWPkDxP/dxz+J4/3ZzCaFvVqRegbhyZ2tzEI2pH7cIjlnCv6HZ4er5A3Jopet
Wz5a31g2JBMNt1GEdxKqekGkWa4eN90G3aTGaPi+uU3ntxR1FzneYMhfmvODAkoE
HIdITTC75LCQICTOO7HLV02+IcZ4DcBogzMc9Z3T6U2gM4pU7L3yoGOvR9jF/2Ct
jA+YDXDT2C+DK6ficX7oFO1i163VIJPe2U0lzSJubMxDlQiKf9grZUlylyQYB6xy
pjmbBVb/hOgEA7HF/YDp7tPmzLxqh/YL1YEOHwsnlPF1eypK/sDtVKhXeWmlDTFj
pjB7VHAe6hh4S6Zwsl9ZxNP4or9fC9BwLAoNfuQQbir6gIloH/Y5SfpcdKsoIlkd
N/w5uajRqbVeESChBP3kQ+iPmKizNqUQscnHh6PK/kM70GEreqxy4pnxodVFTme/
+1NF73Fm5BdINe3QKOhGhkCzYyrLXoiJiHbzqZjJDTkhMfSHVLwsYiUHTPwYFuD7
WAInsz46iVFc2MmrAm6aH/TWqRs/UVIsQpIgKR0lwme2DcF03dUkekWydH99tMLL
bn592O2MJnhQVzCyInu4jhDFi5SmJlb8eOumutEr36+EbVY65m5N7ymOPiotiRwh
k1KXx/w9BxOXOR743fpOazaZkFZeeQ+7QmHS/C8qjKa8MqghOZOrHZ5HbWpE/b81
NTavf8EXn+mJtmWelCblypGZNZrHOwnWdwT3urnelx+b6sLl/7IG4xxczm2ZzsKB
+iO3VsRYykHjNBpMS+jYl7QW91wzbvgbkNqeq/2EEL4WYk59/rsyjp9WlvFGAXKY
ivO0BGFd0mUkEe2INOAxehUlLmJ7XhsmJWkEvZwt3St87F6D8h52bAcY3xv+PSnR
0HpHzsudZOSJvpMvIEZnepeyNnPXBPuyvS/Rd9K3+v+SNwTRILzGvPjxEzT8ILo1
nLYQ58iZwZhZRuABG0ZatH7MD6G8vlKfSmEn1JfWWfVECvGutGZLI3gnJqpR31Uj
F0VOtYn1pQVXFYDdC/eevCllw2w85cOHR8m4E8xKbmpJ1rbk80QqRws6KjG0G5+4
lv6ch6YF5aj5U5Cxha9X7LG+H8Mg4oyBrNxKpQQjMzHnA6MXjfbH59R+nQL6sVfx
lADV+bk2WD+UOn5gg98d+bJuC7uIjVqF5J66P3OqNvi32A2OF8d6VbWq25GbCQVo
SClkCgBfySzsSIhCCkYxbsrqZ90kGX0nSeR3xYLNUII7JCTT0aIMSPxEF/b8+YNh
dAMN3CdbeXGpzjGcseyEZ8W3cmFM6yi9JoqRYJXyLk/QIPs2JcTrZAJEjvNacLc8
pyzxLX92mp9gA+bHQ50fK7PQUioIal29k0lx9KsHWvupo5C2SDP1Ri1wiT/CXf4M
qfTx29lM4loL1tI5ZvopXs2K1VkzRI1NwTqYtYzm0HPAdhwGmJdhZ1URKejd08n0
emGkgTrTeW/PdShBlMrY38Z3cfRHYEPskGbAR9GHL9o+SzQcS5eR7tdEg1hqU4HN
i5O8nJwe4MZMtTBJXPFARlYPSRktci2s+sJwOjqZqwPQ9OhS4juvYXHS7CA49SFp
qOVIZrxt3XLzG4+WvqmCTetcWxOdEYX8ydtJXr+HLRyJPWkDcN8HG+msG/CWsSqz
S8sbFBP3QxonxzJHmU3T/XGJN4xZ8zkhWoQmiRcM538C/y/FOY4nNQA7CFkw6ew8
GgHE2uUHSuuk+bi0M/lH2jNwWae5aGGylN8V7AtGiFm8NI5BE6XTf80I0v/e6d6x
knoTjfVnyhfIxJ0zGlNuNQno+xQxQXZiHrTrMy8FwHGT5oL9VtQvtQaQaVabu50R
/EAUY7xxYn3Q0vYI5WunJpnGOeNEfrxCGAOCFPfuWDZCpPA6ZZ4HtPYHY6a1bimA
RjhxTdMewirbQborSfpYUmPHprKyEmkRcYAktDNGT5CvcFhjMrKIx8BZOO0qPnxh
ahzf6X/kPSKpIWJ7wULpSYZP1IEcl1Fmr8t8DENEnsQpg8inLFsTkUWMt/WJbKIf
DrNbdjJf1EEzRCMnQD+3XXa+p7Moi59ICT3nK9HDYm/ixI6VWU+EsXEo6PZ7rWXC
eHv2+SRdG7jO4aTJP5RFbpSkp5X5/VIezJ3jtskDRshxfzJ3/VRg/tuSyGwWbRoJ
Okt9xU26UW4+tMW6QEFx9A3x5r5MzKo+j5HaK7JrJTsVIXUKEiHDjKuP3j3L0oxZ
ZoVEDLJGEiYiaIkYqBL57+86DEXlkOm16ja4DyXOH1/iXF1GUuIYoBZJuz+yhdjg
S0OSKNJ7vRxz7gAdft4coMB16i3stahGIwjY3ndOqmNOk39xIb0oK3VtZ0oXGjIS
JS8Uy7ZTY5bXNr/00qqvH7V+TNrFxNa4Ce56LFHvtNV/B5qy3D0ko/ReOfMuVYD9
u3DSYJs0o6rz8NF/R5OD7MOs4HcmoTh8lBo247QtggzsDws9n6jwePJyK6mb1zrp
YTkWdj1tQXM+TIEHvuvzj1hjL7WI3PZUottKtqF4hfEUe/tbVty4ZuueeahMTiDt
5A3nljGvhYs3hm9qoqiDUF6Ab7KsfeLR/xRCr6QueGZAbaHEyqG1JFqJi5h9gZol
UEBc6hCDXp8ROP0CPgO0HNVf7ZvbMOPKwnQq8qjrBSJQMTYIojpR/X+/EG/P0dUE
0n0BBrsAvzZ+czRCXJUQIPJMv380bxvDefb2ZnR94wzypLkIBI6ohZhhmFgbAYH/
b0+nJQHuUuaYJ9Az4rtD3zGceWCVC5fnrl7TdGmAQ6VMyNiidn5W6mWXFVu1/rxp
zAl0joOiBkZ6H1OEsMwyy8v4UQ1UBDBank4WE3u6XB/xrkUCE8UiUuE/OTeVUOzW
1ai6Zzd7D64abQklxdQv5jIKiytxta4nca7qtShH1a2wRL70+fowapphp7Rr/cEz
hFkyVW1F1eYJOj+VhNTFjhj9vfMEsgEQ/vJ+VW2XBfHDtmDVEXJPv1tJdugxbMgO
IzcRWtY/leQLAYnyaiNAKV/MvifmkYNUvJ0ZIuZzolno3gNS/Vm74d6yUMQT0u0x
I0uohO2h5IcK1AfKTf/90AFAgPPLUMQXeHhgzZxp8OX0UTawxtWP0D8OEkOVJiE5
E6rgB2FIhElfAZW+KktuQrCp0pjdK6dWaHQBEcDpyxrfVvUIFZ0xBP+A3nwA3xaO
rC2l6fNf2WuhN0jJVQZrksnPw7TUKO/pOoEdkDzX7MfklcGLfB3G1aIAyp20pP6U
qqdn8DZK89YD3tPV7wH7JhRUUhZCrVc7NxcrkuHpqKOdsO7KKModnrurfxbi4c3n
B5sHrnp3P3a3jNe6TvMYgQegtWMKbHzwCtF+vTkFMG3Sx57Ogwp9Vla6/p8SRDpH
tpTFJmMoT0pXmfBCKO2uXG3uetlQXzMv7X6B4ybzsUf+Ff0ljUuz3oqF62eZRBTI
cG2r/c2crNM6zNk8BwfZZmHXySvktHzwsQryqdT2QY2xK33yj9ipl21okl6W9YgG
RG/GO95mBU8fTLKV6wGWjDMBQ9Km0TnnPtzJwqWZg5g5uAadS//863wVFVzFByfC
eIdmXtw2y4yaZGw8jhUKAA1vxNIzHIAb45iHalmJM/8pwaImxCqBVEseCzXc5IKX
i8D/a749UxZDwYiyignhRb2wmwoY0SlTKpoTwX4lka5OmgvD5OxX9hwhI3aXAOdN
m4NTjPw66AAFJ5LEOy94XjwMurMNWh6JV9eARbdqozzs3fP5lkw3Em69ZMlqDANS
ORrALXyr5cGdBJCo6VENTcBOSu408QzP4Mhly19KLs2zFO7k1NMmpSVAMAwynoC2
GmOOnkaSJT5uyC0Yb3HZ+hYJ8i13FiXN35Zxz+36L1pkJdWHk4BqPis1w+6SPbKB
ysUa1Y97fkmUIMj6daj/wTBCptS47yNQRcY2Yps8slwehzyM6tR2Wfyd69h3ndMk
daLfrJEG5pg7uLEZCxK0kH3hiE7TVmjZ2Pcm3jwPLIzD0V64qKLntpm2nW5OdCVv
S8Qi/vn144v9as9nbMtEUaomZuDXjgXzzpKmkAblXyFhSw8LuqoAXM1H8hL8a4OJ
vSe0J7nzc6oL8vkEJ/eeR0w+mqAjryaZKttvzRa/1EOMTGJ75YQNtjK9vR/aD7GJ
1su6++nGaZetrZMNNbqzV3lZU1+8y2XYLX7v4KAJf6wpQwcOtCL27MCEJ/T3r/hN
FM2XNTUynDzDX9QWmXFxblMj2Qooij2eKGXRsYQmPwMEetrgP23jqdwtQ7EJNFGk
c1rytScDLaj2NQqc4WMk1djhIWi+iLxw9choj9M5qT4sEObXINCxj5ESx3aHeOl+
ZfpigsUAj2rhFff148PSXp97UuA53aVg/5L5DFDfbhS2uZmG+lo1ZFuIJ7DHSQdV
zGpVVdLtd4+U2cleQUCY9iFDxNou44c46ILg06RJ1khi+Rp6prKWqQatzS6+CNLr
Ujx3lX5bnkve0flf42xOOBb6Z1r+LZYpmRPGxHui8uTXdzq45H92IK5HoM3WDfrI
0fV0pQBU1xPuWmrhCWaztZ6MyG+jApAFPF48mnUseMjNywtyq7fnWn4LR58k9G+L
GMgio57yNb2e6kpc1x45kY1gZ1GkUl5mGoqURzmHl94efNA8l+AA64+isOyVkwKI
QChZaYPXtFK/rrEKqNFBgO+UWugxq5zbP63vFk2IBiN2M51DezSGj0vya4Xs4AgH
vRTOA7wzkxseGx6fbQdydw7p8XJjx8BeYfFIl9tmqspPWBcMiNlc0hpUDEXOlzYZ
dcyeJX0H84l13FnkFBDK8q/4/uVNhTTBbYUwxuu3BHkcxibkNqqjOKqJZMaPJaNT
65A0lynclDZvgNp1GiqFRxfQlYnkUfvPaAzZLBmokW9zPfJbTO8IT8WVMf299yH0
rQbKUWPOyM3MYKHikUfxtCMdamS4HUuwTQ4UVcwCE7Ae8uiWPSfPh7sLXdL/V7Gn
7qDmZ13rtyZKQPFWU4pUA7N4TLAQH39NL3UtxY4jEp4zv4iOlfLc6xXOtmS1s8j4
xgNpJ5H1z+02abG3MMYH3zyoI3/wSxzW9p5o5VZVAgbwlfhnGqGzJ8QQ5KyTUBOc
ekQldDt3gMn6DcuVfxhQWKWOGU/Rhp//9DE6p6aNJnNyGUtXnAcFMmdkpOkVR2U1
j+O/Nb9Qe/RRrwl4x89J1b7o5QE838fv1yugeWELKA7lH3B0GyvVlEVsog199Jq7
POXIum2Q4R0GXPzy7GrkktsVMp2syeBC7ef+eyhug++YM+lO9T+mJzpmFrr0CzxO
FnE/buWN8Q/QnLohMD4PloSvOcc9RLR3HspoHC6UyEdkGZWtvuKxd5SYzE3rrC3O
bIeWAZYd556St+WUJi0NPCWSinDtRerRT0rZn0Us/nya40Gm2tyXLkuJwU70zGYy
qLsCpJSFS0o+hh89B6iVS1FKm+++mGrg0IztxfRbptxFnD0LCzr8zq44lFrvI2Jv
nH0WFLDssA9epRByHzl5Ma0C+TIhh2IS1ruEcykCny3zV50GIe1EvDuhEzfItohw
5OJ04nxFttrq4IinCpmv8BmBtDILTRB+9A1NqQV7Y2n6wosou6+YKzLBxqDhVJqh
+n92XcZsYmpEqjF96UVvwFSXCFrNKCcjs8JDBRa79dK6+XOAFizPZmdF1XVNHYTi
PEz4El/Iu1Ukf1IBXt0ELrmNXXLIv862Ym0T82fVLILxAQjjt1cW4/RZM3iFEG9Z
Em4jrttqo9SVm1eV3urPlkZW3A6eBBTbM0OgdFjLM/D5+EAiRJm9Ty2IYFStRw8w
P44RZwV9gK16vssrsVanOz10qXat0J5t13/eKfkIZ0GQYQJ1M+4cSH7p/6Rdggmu
TLxeFoedSm/eVSEzTceOuDBV8cteujDkrqWpz87kiohQyaY6BqJgg0RIXLRwogi7
38cDzJJXG+Th2nKTypSSHB0C45f/1t1Vpz4p82MKalUaPGo/576PYpW1YdUbMh7O
SMWcodFPUOAtQRWUx3HT3HPnvqJdDs2s3v5Ipk1xFtolbZYw0VwUo9v9nQrOO/do
opVyGVEKWrPejiX1xtPdRN9MdEw9udRmToYy883Q9FHNhu3WRGeetrfO1F1Y1XyF
GxmImfs+Md6jcvPehG23Dq7IOJ15FCjSH4tapI0wXDW2b60F4TPxi8Ko3ADZ40XH
CxtoNqvmPG7nmeCYKB4QXwtz14qJk2OLeY89dkwU7sKPpXfv1ZjD7LvcbErGZGAd
1i7hI/ATqNdLbNm5wEkxjO/IfUeIR1uzp6PMqCxEMema51EhPZ+0mQSKbb+Z0NxY
R7gFuoTg6QCLdOGqu/6CwWSuTV5eh07n4cP+uhqcxTWT7Wb3jBIwRg/PZB+2U8op
pJjxnGQGsjivQY0E/jx9QoS7TjekAEobm/PI6e3c7lu37K8CeeJtJhDrUoL/PCB9
fzAv8clZjHPnCVqfnNo1xgproB/X7zqTtvf8R/VEgIwvrkYWvx+3hVd2hA8QlsCK
zono3R0U4DuPThgSWpDA19x7rH/RYN1+ULw9Wg4Is7qJ8S2Tr4xr8RtRY6mJuSwL
n0ZZny/6yU/P+2VcIf2N8exPLz7JTRqZ1sdXlQuah0Ktq99XzsQEH1xNgpduD/Un
kSDAFZN5eAY4UDu5z+qVK5euKOkRKifVQ2IlJya56B7y3JO6jjhmKE1Zh6jNWk3V
U4HUXzFf732DLvW3MMRe2oyXMeJWqYHSGzaIBbaGLDrjSEFLZg2QYeSXRzC3hfwU
I/iYrUzYmi6KI4d8nWmgip1pd3olv80GMd77xVpmB9M0byw9rHs1nk/hAsABRFGu
OUBQOUGR4vt/rtiJL5J7nEAsgyxPzh6cK6BE69E4/mksjWChoIPeOdmADsXBmHoN
zyhYOBqAGAmvE+/mm3xrVsiuUIarzN+7H6sMyBamm495tn8Dnoyv87lqYm3dTI0H
O6Wa+sE18NeTWZbROLJgfTAIYLcWmmlx1EZADemucf18Az5Bf47D8y8ijhW9CvuL
XXBiwTkIavEZgEjL+pm0aHOONMUHfUu9B1e9Lvxv/WxYd2x528p1psjuDe1/HrQb
uTyZlaowp7p0iC0awFRv2qYk04zgNtdEzAn1ngiDt8iiv0cMUv8LiPQAy0HcIZGP
fe7Jh225KjCQDymsP5trHqFzjrGlke6z8hp4JELKprSU86xzLt61/1k9ajXa95pZ
P0YeE7R3BxUXTqfOS8SEgZg7NLzkm6sGgRwC0JdJeDD4pgeDpN42LDu5QJVUSED9
El56oDRO4F7SpIpwoccVYdwHbn3nxgA3gUumj6EFQMWgal2QDbHTNbwvHK156/oZ
QUy5mpsj6FQemSo3JVbDdfraYmHXQmghlIKHczM0H/Zp5YPKSWL05ZFpDeNhko8A
+n+AECksn8q9fUojcBBOmYGbOwhREcrN0sWhF7NhaA0ezFp8dBDebHxv4fqJgfqX
F6FRKFgv3IQXCGMhQaimMFLDWZGMOYRDB21YiY1s9HXWKQDU+yKJcd+TWlondmJe
In567z5UYy5ub2rfvIhwxr+GhUtdcKQIdwppLn4T6PR3NA6R/0DjaDwF0Hp/mIa1
OqAhHFiy4CidU7IFFKmEQIEEOrqoqQsygbFp0m2sbCZWwRyskEOGk7fvSnOIL0Xn
jEFatAMvagPGguLB4ZnlsSPJNNornDNrauwQEi1aF4gVrlOtYKMH/Ghtte3BWzzF
2G909EPf7ztqeYJF2eXUOJw6FWhCPw+fnxuTKbuPNqtm1KEmPVKhwYa1Jymg8tw0
xQQ6XkhSid2b7IqzeRDYQOKYH9Yse0hkUjgJ71jGMQA+crvKLjKbsaINOqsJwKRF
UXKznH7eZAQ8klnQU1cXBY9jjEiwIjpW95pUpNWfuXjV6dFejBSV3LyI1HFMBTKj
HQHxMFFo26JeAkcse7xt/8j5LpxCisJvwXPgJhrl7y7ngzIOsteaefRMHDKyym+B
YvBWt5NCvbJuuszVchndGGAV9qayesw3NIBYgbIH/KMs4jtJRoZkdu1NuPedBiEd
PK4humWkiuMwtWsLaTZGnJ5+j+rh+y9uxVUF3IKcs7rEs8YlTunPbyU4r3aS9WrL
o3mmjsvXWu1xh7yjZFONdoAY+m5a34vulA4QHMxS7n1UdKcsrV3zkklxVXjaKlTa
Hqb8TTAFTlVidiUII75aKzXcANfhLq5WQrV5tc6SxngEeW4TOKuw5wkuaVEgUoEi
dhF3gzOWjyoEXGu+MiAIjPJDtYeIcU5G8uGxfS/pU1vJjlTKLSZ+PgTG9gYbDmF2
BiNhsNdBGkc7U+Qaa+PnmdA66AVgVSHd4lmzRgC57fCw/4x+Qtv9XRltDW6PknZF
uTHgu7NuV7WXxYQXsfLf69OXOramvcYVpevl3AoSyE3gDK1vF3ejnzHXQGSTAJzA
NtcqJvJ8kVnWtbAciRDIQnCgS1GoBT2dVGreRY2StcKylr2Ae7pl21bkzAZzXXya
WwmmDZ4vXwDU70mqcHVvEpWSEPB8tw3AzIKsyHoTnErBEUOdG0Z6XtiJ7EZQOfOK
3b1iwVAxK6aCSFc/3xoxvptGoHtvFsBLcyTqukf4sP7foqPgW19ZbVyqtQsNHw/1
Y2rPSsMTqujZCL/xIqJ45iMZud2U+3CNeLuh0Q1XpYszAw+c/Re8M1jwZrVqM/tJ
fHMFPy2f6SHlbd6FXcONcDFv2RDnpRv1fAQNWS0RbIK2NqjtwOJ5NkXafbVdAKSA
hqrdPL5dpO7OpDK9YbC8OXOxQhnrBxmXCl8HhJBSUWfrGw62KuCk+8oo0wFtuiEw
uR4jKWRrmfgELfyhC45mB8FUidZq97xAPzrVauaiuBbhbaD3gk5Loom81+HSnbfU
jPzuXi4NJba3vfxuKEmrLAcVavAlgoXWvR6pE5zBH3sHzUALrxQYMtfXtOc0v2lT
eGHLhxGOGsPQtI2LTwg8p4mh6r5a5Njs5el4+Tyk0dxhJKhkQEcI3W4HEZzVKPKF
M7rzo7njlZPbxwaXZLT+dsEs5AAJrUhV+N0GFXusPzd5FyP0Lo2Z+iQlxqZDZAEd
QJN3eeeKiepS7nRXh9SdYbIqOESF8CJ62TLldY83Vven1fZCFJJNB/ndk6G6QjBF
IiiEUwDG33TYxWOxAK+/RUsW6dlWwABN8ZHXLBaxPjC5RPFUvkXyw8egBblecujE
vWWWPwqClECDEUc7zP2nfSqbztQUr8x4js7shSSvrpZdK6Ns5rRzWmlk+OIPAeWZ
G8voPZMaPJryBgDUFwrIwoMGaO3sSveIqp+fEr7oRQEnFIeAnnC4BLQSB9im1DI5
IGgEKFALuxgjG2c4xyUTZlrwdrGLSryA1XGHAR8EBybofWstR0tF0sAjZkhv/FxL
VGc+ShHl+U8y3DQUOzuK+zUevrz4BvtrK9k8/XXw3RWzuZli0LdPpS/Iu/7818K2
F5pRXLmzuyqlCaV1HDhMpcwVZpF9y5ITMjWeltz6OC6+1wBLlurf1EwdBKYY0jfQ
td2YYF3pWOtctSJyJiuazXgpAWVgGjKXeRCiu2UZYEovbZc0Q0yitwgexpmT8siJ
Wq9MlDpfpY1p+l7LZaGBGK32uLMmDjmj36ZsDK7yAol+XD1zz8MZMjnB4odfwdof
s05rVkok4pWyvx9YdTck8l/UyiJbbS6kbJgy48CKw+dXAoY0HRO7nfulYcZuuCg9
toh9At3ZF5FpVjD9o4QoRrl7cEPUsrlsqBq9IkUx3kh16MSDdwfniej1aTG/YgnU
GfV6yY/9ANIcXc3/MiApkOYEqTA06hBXm+A+O6JB/5gaBKmXs8MSasrPOzPY99fU
Kg0T7BPtuRhMhHohMd5f8pgxMKRxjSpNZD3xUWV4k7DbyvNOiVaQivp+np5wwuvY
34teSzJ7MICwuJnBPIqXauTpXWiA8RXmXbTSxt2+W/DOTVXPZiDuZxG3geE2ioPY
TBQPYQ1QInNCTek9EW4yvQ/xXo0T5MCDB9MD/sbVqWfwTrx1nourqOo/7dnM5QVS
w4mX3S3XPm9C1Hx6YzUNwiL39ryjpf0TA5qySTJs6Y6UKhExi/dhHLVv6NSW5869
5qgAmBWomlGglEF9Y/EXc8g9pyNUNQT/vyhkfcWPFWm9mpjFMdAkFMaJOPKtY3md
lL1NO5tXJlNWOBQpHNO54ANG1jiXxhioklvA9q0LOYwd7Uglm0+MssElQtev35Oh
BvZwq5VmZlUTQyS5qycjBQnHNRt+PwXaZh0BdL5kj7g+NW/a0jEJFhxOyk5XqljL
qFw2tLKG45to824gYvaIXoXFSON40W1A4635+kCbm7vcrTzsNXyotFTvBzuePPEY
747LfktHBe1+5UONRwDXgqdcP7tYQB+n/DHmlU0k3YnXXl7ihsDFLD8/t+6riufS
l6f0IMsFJ+alZzqNSgX8zxLUIrbyf3jDztPP8nw2pqsyzbIJmMEZfpg1lmtzZfwa
dfocPCiLL+geQhU3jCOFBo2Y+AH4e/oH1qhzCo2KvpDORa7VToLxUYaitkyuAh11
alA3bHdkTA5PufnEB5zJSD+ZprVKyxq8onwUbY8bERL2B+1aSGbedsuBZZgeTXA+
gYYshBmHrZyvJQXXO4xly0k2AkaJWUoEo9Mo0dFlZZk1wOwuJTCIkrx4yZn//keA
nZFElyqloEn+Fj2KFD2DTEJFhsxx1z3AjAh/jS8QuUPmEfKqChJSfnoDfyry3N/R
YbTNoVGul3AaJw1swrxlP2TP3dNx83kvqCkuvEnTFKFroBZlxWygMSPtGpyd80J9
rZqZ39Uxw5IXaYBO9oZO38HgGcJ3hHtOC8xv/94sA8bNEtK+CB3OWRYJJ8jJ1GaT
Sy7YKig2Krbrm+ghhOCA+eJzruU9k4cpw3yZKph6XPkYlja9n4SWOWMzaufVCObu
w77lfEh+PCKJauSC4NkC2SaGgdT2+A0Gh0t7oa+pUxVt4jq2/AghTkB2yMgJGgGD
b0lGGZy0cUozpHn3YX8IedGA2tBUA29ZPGkfjF4KubrNtJD6UKfIey+1mx5ykUtX
pUo2pGoSTnwvvzFA9DmU241St3/XO32eVIAnnFzh6iD0qnGNsOpzbAb43+0+06EW
6kFvb7x5yP9R99JE6a04bqve0vlUmscCayejpDPoF/2NoBZ+hNCaDyXZ6Vnb1FLd
CphUX6Pn2nAzHkiSxV2AkS6Vep9zWfN45JndVLb93x4zQOBecYO/fTIxIsHGHMx+
6WWnu5oGrBURlX+57coeW5VIR6ehYvRT1VQBYW2rErvlmZg0RWxMy4UN4SMCWRDi
ceRhD/ODOILo2Din1YHZVeLLguVNlqpNYaPhDvH+rpJKBux6H4c29iNR8M7gIlav
E2ZzE25T8n6kECYqS2lLEt0D4F6xb6mPzX52oP00IVa1kkLupFEt+TnRxvOhdVBk
4Qfxq2JN0G4HLn4Zr/R46zpJzyFNZy6yYUrs9zA9Cpu7302Tkl7wFOSzeZX9l9QZ
Idew9+NrZj8aaTb98pCalS9d4ydFDrp48xB8je2kapbl1ANWUwx9/LmmAZH5LIZR
CHB6s1GdK+HyFrf3Mk7TlOvoK35XM2OZSItphc6yiKXjgbI/grqbCrjgRt6vVgF+
QFNY8WgaXR385yt47hsP6RUy9U7xAeodgXc/nbBMxnnnyDpF3WM/kk9X+3LeUDF9
5mHm1KEK48TVrB8lCB/AwohDuXiqqNMNrmZlhwUux2Pvx4CDfik795ofd7lCktO6
Fwrr1lRqtjL56qjwRHh1psj9+U3WtDmNcxhDMRAQHcFzmEQjxTjzKahL87oY/oIY
SBhxAUKL7K3BMiZg65exPdpvrp430IXk0pe05dgWVYVZmzMRrvm+9bCOZb+cMp1O
/W3dzIi0Col5Zf/XpgW+Cs5XhNm1l4lj7ZyHO970zwiIYw2pFF3YhiiEhRPOYxPT
ai0tVX04e1D5/4NmSO/dQg5W3oT3Yj+vRmwrNCUi+C1hUGh/oI4cXOrnuRcRObWP
p+t57AKgstwRYHSCTwq510/D0jjm2if/8JojLnTpi5o5kvbVrTF0c+6/wSaqgROE
ImzwGPwgACYJO8Ull3uGwq3QPrP6KATyh5Rm7SPBoZ/rzduSnhhLcoraczS1MztE
pTlv0oOqUZJ8NxFtMeN8VX7K695Te//5FEY9R9ElZ2kDmIatMZL74/WFkIDUBNgk
l1JZ4/+5EEH35//9tvbNENQlIJ/8N6qBKFXQQDpOR0QxK+ZJg9WWw4itNnz72IQK
FAHs+v806NdGy11T5lJLLOweMdpQj6/B/No47nlel0UMWcHSrKYfh6uaRucvjH8X
8JgG6OvxucLW0qJ3o5vGPHbWPju0rYDIOuwZljj/x6KlSNjU4wALeKWU9YwHF4eM
FpQ/rSpOGBzmR6OBB7aksUEVtM5kX+sPxsspeY8DkhvZSzoTcsu5wtwVBeX6Hko0
tnXRmXyfJCvN0izJN3ZIDqq5RzjLgit/+2qhT3wIfaOxKs9opP9J54dq3cNkCYth
v9OrNCSo9qw8L0ePyi02lfpbg6ZRcQFhxkqOPc4W23wqKRJCepTdlGLbHnP85eUq
O2BnaiTwhTpDmmIbnEYQgDV2joS2gfjnQR+A5im6OYRpWjYXo0RvFUYlI+9XZf47
E07mVKPNUbz1Iczwu9VqhQZKY+EXdi580G9m+Y9gTZam+1jdlnoCovwpN+L6uMWh
4RwWT0qV60ZrZeP/vILhPofP1uTDyUCdWTsxPPMMrRd8Bkun1at8H/ThC5iyMyVs
w+IJwG/uYq7gNHVkOGk2R7/pV2knkMyCVuHEyBKfmS6nLI16p/VsL7eHVaJ4b4rh
EwbtPmmZ0F6fkyuD5fQcglVSv6r2Ommz1j79TEIzEtWoMgvsY+uHWFxDC5S94mnT
tBrrOzvYLhkkMk0qfv4W/k0cq0r4EZbeFbFSfEg9r68gDXnT79fcNcvNmwPufUyl
U6th7VEWDdfqNSeKBigthmkZ5MBFxnBu5GGn9ZpeWW+hRKvIUt7cKhGP360Y+vcg
cV9UJKizi2BvtvfuEoWPic28gw7xxev70EsSdfATAXeHAkNDXMNHAQWQ2pj/uGUy
Tt8Gt8/lvnYlZhqxUi71/zphkJMfDYNQcH0AWx3dtHg+1F18DNRlzbPgj25WE6Uv
qVN4LsSZahRxBZqjsRhzR3k67+GyOdqsEMoBmg8r7s/7CvBSxm7riw/8uFxV57ss
M+dcSkX6Y9Mh+SrvjnqlUoOWxPIX491XAH6ROXrYWRPLiA1Jv2Kwxzg2256gDPYm
FRuYwIKev30BQWbNHrpRY9p/Ii4941A0ymvw1s5C6zYsZViBX5jgmAzlWq3Fa3++
jzNdF2lLinMoEdp0eGvI3EJhEgoWKqH1ruH8Tn7CW6GmcLYnSbl6Ybx2UfF7msge
h6vRIv/GsYSIbw3MJL7VFHcnDdoxf73Ehroi7NGFd7/aTw/O4TDY3Cbt0R6hQyZs
2MU1+qbJrD8Lmqalb9hrqcpe+ZXBBUnpjsrcsFCGHxXmi8a8cbCffV7CwGKxIdDv
6NFSIiwOXsBVol8muGfIJRgfSpLoR0+qhaK0Pdvd/Mbze/U7dAxVQlfA9SbtFpm4
ozizmKuZKIf4a5N+Gzt4YXdruxcADX2qtlFB+Y7TWY5xKqoKCkpgMNaXacodF1KA
aEqiVfCIjNhQFDIXJGiJuN+GMUuFTGGlHDFqumT4OtoBbDdr+4b6zw5RCOArGtiU
MQW0EMnQjDtX7AMz/jLaUSHgAfMfPKU6lKL+fJT9uhKFXDTOobIawxxO6I8+690k
IvHpyPxnQ5Lxt17EkkfKHIPyVsirR6BlqfZ4h57igIs3itNMZpPXb5l5ycL/GpxW
bWC2DJC+4FnGs76JKlqthFBxEZj0Pp3dWR1xIUE3u49LHImVsdXuSz2YOByrzPzh
SXxuTii5WaroB3sYbmdU7h0Y+/77FSmOq1RNIhjD2LS9lSiFDXBMReaHmad71i8j
kYDOpqSRRc8DzPC/5Y9Nc5XvpMdwHp9oPkHXsGqUWQnVxWANqGrOK7Et+coQMP6u
XW6kxu6Fmj+6WA10lihgtAgLECZrPZYdF0o9b3dOZMaATbdPvIuXtkT4d1Q5jtvy
ItvZ/mAzTU2Q9G4WL4JC9QE1U4pe1edrGhGnnc392Ig3NS6aQjRbXneecokhFJN4
MBolzpHD/tuybR639h3Md3OFlxCXv9w6jRDaFpuk3C6F9WswKhbeuTkt7REEhOok
rmk6NfjIwFaHDGdOIPWf+wm/DgUIQhSWKBepfbVnWZ6l6XZ4QW9IyFiu1zwO4io3
3SbyhTWk8tFTjzLZmOEevUHCjohHaGldJp8auXM2e7m+ZRDb/ff4n4aemxr1uQvl
7u95f1FZjRpY83z4rexuzAXVE8OZOXpWxQeXA9rfYQXz70A7F8SjxV+YMGv+o/bN
B15oY2ydTIIH/77/tSYyioMH0DGJksXldupw440RbojwLQE76+1GnjgF/h/Oyvqk
OP5e49HpnfqliG9EVwTeOoOszYArshME1QD1tIQzTYrgK6Ywmoo5dgrEgkqHHLH8
Xu7oDwke+1Yl4U5X+38orhMu0bayh3XYLeYEQ9NflFXPrrsvC6LX8vxeImj6UWFW
LfEXwgLwsMODmimrLcW1/hXjB0au+5+XnLVlu/IAmC2oOiAdcBwViHTFv09MqqAi
jSTu6NONsZi3wxqIIOYsk0FBmgkrJze9t2laD9cvwFcszEe8olJeubBVl4eSiGy5
SHrPpWbfupHARv3mnmvgvRKyr+ZDUnSR0HQoD3GsxQuKB+Zu55z/ahluL8BqbZRu
acKgMBA02FKGvKaP9j805QrDa0H8+Ep8yPGftZLzpjdE8Ii5Dv64cV4jQ6GNrhnW
Vsg8MgjvJLMlGZQ0NcBdLFnJf2Vh8V4XPjJhyjL1NA4wu+IOz/PC3/+ZxGnWw+bq
Dj4KWyNnqeZHI5zoi5i1pRVpqnhf3lsjvAtQ0vFfWDu7EvE4+23V6De1qSdNSYvL
Q2yVlNZfi6TStc6YIjJjtDo4ZP+Ms+diBif8ZOsA/4J8eGl3uUE8dSXi8taU6lED
TxPiXnOpNyvxYqxvL1GOXBtmK9cVOxfq9qedrCMCEK6eSKQLohVS4iPdq2cOr0Fi
ukJ8A/wD83fwZFo8eXYDCueGjghZ4mm31vNKCzLLe++oKXP8xuasFthXirWFxRab
W+2DN880CHJCElqnBrKGzYFuHscFCi1ujW8gMkGeXZBVpT2JYyedEWZZc0pKgGKM
k9V9ys0SK30UJ4MiNj6ryhFKS4gxTDh7xySUsEJCPUkQevtUJscJFJT0tGbwiq2P
YWp16fH8DKkXPNFSVwg+2oBF9k4djiC7B4oU3tkjhEaN+H1XfQO/79TrluhBgQh8
wfmiN8K7qpE2M+KF668oprmL59C3sqKOwB3rMYCT0/lm6+xUjLo9I/ljjA4HXiIa
ZNdcOGVPXXWZHnIS3bwtQ/DT9UCiODyD6o0Vk+lsnByB8ITcNzfroy7eBP+6TOh3
4AVgrHwD7ijucTFRDzALgvaQTAbZlFg8/z9WCFEJ9Ie8NSkRmafbScxa0U8a3UF9
q/mqr/ltNF3qcKhnar5kyd/WrEoPy67qiEIoQ0aq6ypqOzUT6gbOOQtFZNksGbjz
XHQvzLkDqK8KLQyZqqFQTNQr2rzwBm2niATDLHnlp+VB68O1aV5ewuBiBT+TakeH
idEtZMzUi1sWkv62OgFDifcnbTTm4LFxr3m56LX82RbXYHkQgoRlmwv4VsOK7al7
ewTpJ0wllbs4VXmJbHWTDW1vWlYlGcCvapJdfdLUBHiWfKiI/eFAbA4D9w4He1dD
uPZWkX+CYQePavmh9s4lQBisxqhLj+6TXSVduD/Iw52/XixTLjbWP2zy+isajUf2
fSb2Eryl26MQeNidui7gHk1T3iKkIyCeg63HejvwS6ewUq5H1eR9hl+kYpG9lq9j
hqU0Waf9bfezTRq8uVIcwfmiQlKtBptYqMOIX3SLYPDUZbDF1RGbhuUYZHMdSDLP
BaL8DfgDMOpVaYbUIttMW909q2/3pxCnVgclZbeoSxsWdNu7g06puV8V4JOZdwjp
CXSePx2riG2zvLVtR6/vX4Rg73Y7jjichPzX9A9AiDEdXQ49w+raMr96GAvQ3z/2
TuZKLFM29wrEyILtvm0oUdjqh2E3GosACwOrq8SKKK8ppsduF2xXtMMzhd/2CO2m
pTpCAo5MLHIwmtCJJ0T63whr7VhLZgONogH1cCIb76Tfbe3KINMTXcJioyHjw9F2
jD1y1hIMOKNgxgK/hc2iyO4ZK+QsfewXqBkienLt041z4rE5Ko5VbKgYrwbxaP4U
9Heqpcjq4ETT0D0QSQGYe3FZorF3XAzVsbqUTNoa6NHKsh6r49jdC4sSrc0sQhah
H/ifBOD7/ebXFiA9GV5wQmAoWjsQJQ+jKPnR6jQQ1sBQR2Yal/PtrbeDTjeiz84j
Re/FVkDxE2bEn5xttDhuZzfkM8yzJLWfiMZMz5DoNfCwFw/ii6+Ijk8bhy5kHIPq
W4fYIESCz5ZsovVVOaCSMvbwLztvYVPKUYeBKgMN7UoyuumKGpUwG0b6XJVJ7ooq
tbAGkY48ANsrISDAIf8MB/eAUqhIDoAahl71Uz3VEuXN4TghCN70GkLHQ5KYlZUO
gPFEJcdv//T3/pkFdxWuTvgi2rt58lqCz8gkW5x0+bbjaoNnAgfjjO29SKKRMVKK
GiFOGV+lDL9a0A8hpVoBf3uu20lp5UWNmUyRnaEwuPrAbjWKMuKWhxOzSvAqoRTj
QSi7irtpahjsRx90D+W1IAW1YF4J17ncCMcq7pbPLS/H4tBS9bUMY1YE1c3G9IQv
zxh3548R+IL0TeEZs5NS3SMBJ0YfRfOdAnM9vLmgHmc4EW+5WFKdZsHjAmpZ7hfl
rBqhW3HFN5M6bi5iGQ7RlRlhflmscH25Ee0aD1E2RPlmoy8IHWJm+SkC0sZxXlf4
IGV0cy0kJFinGSGYhA2dFEuWkJPn7R8fAR8FY2/1mzOSz76B5d5WfmPu/Z+C/kxr
qMH3aA/9MVVBj9U5XT4UZvk6v5i17kJR8lDWsx8ug/F1MyiINWSdsVH0FnHwzHSF
B28XAGAzkKQhpoK+W0d6mtqAGYsAdY9JCy2OxB2FjxbHsJMDa4Y/t/6duQHuVdc5
YiC+DI3k9UU3aR1demX0I+MuGqpDy1qV6lqIo4a9NRTk0Nh/EBhou8jpGfANHMr8
Aq6AQ9iklHTmXhtVbAckk/Q3V98lN0QR03FomSklKaC9EXjfB7oqpLBwMMZyo+Lt
rDVf/MU967gwbpr69VB/IuOH98gcBTT+UlcADckrAZlAohwtAkpPuR0GosCI1Fc7
dluBfPSpyZDukK2FtzqLccwUT9tVkTiVJqsvp0urajHXjtBc/PDMT6a425XYSJTW
X9N2pIP+N7kYNWZR8q3Vci1vh2nwcLwTXP+Pwm1WojzN0D6/aDvDF2wqoMaTEDlm
puzMGuOw/XAOtJtcR9miqn6o85goMIgC3tbZxeWsnwkrQfh6Jjr7Y46aTII5hFcq
rLLQ5OQTenorg/Q+yQGlu98QWOLKCy6tTRXPPx0NVlpRs+nx2Iq2vcWupdT3I+Fe
TpSy7Ag6FiP4U9YK8m7zLX3XQxZfTjfXZCJghwvUg2x27yaO4JfR+x96DEHu8+lE
0+ULvZ8eNHj14orJ6Glxu4ZIWe5kYODSrctjexjQJN0gv5y6EzjePmGKWKiN/AeT
joyxlWMehmthp9M+XO54EpINnZMfGGbJ2+C/ZDfq44eTfZIXLofpZqVrN1C2h06e
ltgMkz/OkbaXLbhjzgILwHfyjRFjhLt5PAfcgu6F2Ed6WQE7no2GiM9E+Vi9yVRk
TScX7SD5c6TbpQ/nBsga0reKHmbXzdoakuuox7ceuN3OQz5LOzwOEBIiXfwIlW75
jkNl850aFYlMH0N+B86FM8UKZdmDEFHBuf5MfdJeXFBW7Ro3gtk7npWF997zDOAw
KZJ5BmosgJ01PyA7DJVurWLZ/u/yVHB7eYpDbm+uPZT7ATYZk9IPaGkgEA5t6TIF
DSeaAbLxfpbx9yjbNDHlkLoe0APl2HBdDPZm6nEPprae8cqt6WhJ+yYeZ/zzfbo9
1dL53/FaQuY9dMiVJQCbvInLpuMif2Qcuf82wH95AFFLBAyUPhdOCVTyTn7JkXFo
BFs4AQvVxWue6NKs6Wn2JugkqFfuAqfHG/Psrt8Pz9J6UEZzr5hIQVJ1H6zqCCee
8Ofr05512Mr1rECal17C3rOoKIQQcppBkQ+t4mMbfmszuH7HcrjfmbJA26JJvame
yOsH8mewbqzPisZabQaZqzwreT4MvXeBObgG+GJqowT8RnmpvYbSdGN5YgyXsX37
2rdF9SyC+4Z7VLdNkXITdzUXYGcg41FOO09+MVez+QSITnPSOwtU2/XDDDw/MvbQ
SPK9WwzXzMw/DJV5CoqwMvL8/o7W3X+bYRkzcOLXI4IBBZt3HErjQGkY3kndX7X+
vZuOpI7wmM+fU/NFGXx2cjAkNQJI1gSOCZwrvamem9rFDYupTk6cNPq/t7g3yJbS
qXNZoexriLS7pIkqLxJAYC5fSEKArAu+VCoxGDYiHB6WuplzSEJ1pMwhAWfxu8oI
2Djl53d1C13NOtGzni3A+rbEFAb36aQz+7RBekk/JY2sL7RQNGcJ1gRdqEHwCQMg
hzhW9+ZeMy2gzcQ6f08+Yjoz3cE67kky22rxZxmhZvbcmJv2Ux8gpvcMWoTJOgR1
13SzmtgBgjytkiQ+C1ryIJr78Mk4dJ9pwzZAzuXexeAldphiE4fev1ht6wGoxnur
8Trdw18EJbyzc0/AIhVw0Xp6vPnAkdRfm24hwKMCDI90XA4wINdYQ9UVXkroNYiY
JvU9ZiUE6N61ANNhgvP6okEqVUpiCUqMELamcoXsCbd+ZpC+9YVzoikOCAJHXJDm
4k4ECirsqctTbuLojjQYKSo3lfNV+NvtnbgacEFjJTBhRLQkPeJKcbbO/ndprJ8D
IBf528FV73X1dO4RFrC372k2DA0Ezo7a7J1nGVhubffhTDeuUDtrK5OLU6cglXhl
PRGWQwFfpIOaCjWFNtUHNj5gt9ZpPxklbl9enLZKZXojVgAd9yX7x/V8BD3GwRRq
ImZbLACNDMOHay+eiI2yqG8UOeoAWLeWvTyWYZWoEX6IZxX5DbYocw87pg/t4B6y
IHyuYnj1RWlrHXcMwFJ/Wmk1DMUB0TnfXZLfsH+ElPo3YAZfA5DIvIm5TsWLNI16
vWMRGDchNkGWxFuWJpQRLMRr08g4NdIJxYhZYcLdgVYTnyMUaKKYuYR1MsF5wTdm
ZYOKuOlv+2kebGWON8tStW5OOpeEeeU3zHiC3u0r3S9wrXM+bfeoavRUVYFtKouX
B7Fh8GzCn9wzIyhDDup372/W6PeY/99qPFL8X3OqgIkqytMRlZrRrM3ejNEbWdlJ
WNstY4oyuotvl6rcXDU4OU7UoZ9US5cEg2QPoUHlz4D3dKM2ZuL9odn1WlbswLxM
uu8KGoPbQjI60gc56kBODEYkLlAQeAWvG7ymh9hsMBj2wXB6gCVJvnsQ2arbTCTp
sT2xcsp+MNFGaMhJ8lxUpxTTXdDf3BUgDgzCzT9IxFM5lQx9qDqs8aDj/nb/JqzM
N+ViwuLb9Ff0tAVZOZ4hLnVOxlP/Q5w5izEHj5OuVGeV3ykWzWSw5C5BAqFvJLz8
tiOL/dleX7xOVNmeDJ3P/9S5gq4mow6Q1d3YM/gh+JmCyWn6AbJ3BDnVLjQBUNK3
o7zvTJ74OFfCrOupJ+7RjBEN5EjosSfDkEn2aOKsYw2w5kidFjXp7xB+cmBRY4YN
fNZNwTOSVs1fXUMfM/wKSRoR7AnAV2/0D5rY0CLsgTtxXYqkQ49Xf3U2MQH8E91a
a4lLt6F3WbhkvE0m0OnKsEykOItBcu96tIpEIF9WR+jFF3wH0MQ82GF/U06GAhVt
g7GbjkrHFZTqCznO12pafjxwJQfzZ3gU2npruTK9fTTr1Gha2iT+Qe1VOatqUT+y
viS7a3lFPvdMke2BjPKDVZVBSo4yfWUvsLKKBzkqm4lwlIzjQIIzKb5yR03iDZkH
mYFU1pNbu0nTAn/qCLmER3tLSznD0t/478/aB5F+WCh/2ntKP5P5m7qCsjRXweV2
e60pc++4GVADs5MH5bEtrCbBbThGLNgL5y3VRYOOyeypN3KNPWC5Z3pCrlfJ2qeK
riNkvo+6yMkqz7bn8vIGSHtjJmsa7V9q7u1hRM8qVv54+sVHgS10xtyd97qRrzIi
oPbsbgSC2tceLwC3uEF5qt+NbMRwVVpNpj36GI0q6JV1bQm2aAAEJ4km+sGl8DY4
v6ncGfANbb5OvDaqW/0rGgNri/NjsCd9nx2Kge5Yo29TsMiS3qmGH2NxWnAMX5jr
lBPRMxismXH/OltuhdA5yb2DB5gKPb+j88NSh4TmF+RZY731cX/Bv/7t+YovJZpM
lJns5kkMiJDXRwn7obuoFxfwStRNeh9sTapBJJg9hQqaznrtNCX/k1xQDEoDmgEn
q5fGDBD7H8KSTuooLsLuSG8tLpKuMXVGxFd2pRwCsYajUo4qiudDk+jhwfONc1Cd
/aGOaXP7g0H77z2sm6aeXl0VNeJYUXjZIP7ZeGAdtir7W8lSIvKYUx8DImBLXMmO
XyVsOn7+iBeubDSNZV9b0DpjppmJ22cUymDbXNsrlYcjoVQOE5I43sXGU6OZYsmh
cJ8sULCBEnLKt5MSVuuMw+SGZp+2AEuKAqAVpz3fNWlaXcaZmfylecfGdKNdqYuu
msPq8JzrkBZ6x/hxem9+PS+t9CYK6kfILml6oCL0WtXT8g86N//znUfpH5WFvNPO
kI0IMJH6ZWvAxjecpn7Cic1UAeD8Dcq6zMpIEPZfrxxt94JsZP0NCuTthQlYZQA5
nYXoysL3JfCs/mUZ8Nt1CdGalMUBYLlMPht/xvOpIy8Vs1U+GYa1IjRbIMwZ55LJ
AaTS0vkDFvUzdrv7V6gDyk4hO/bmwxPOSIxFtTRzH7gj9Ukz5ud6taE2S2lTCjVs
xZl9U3HsmQHs3Csy9WOkbBTVY3HKHxfEloeIQLL8V1L5aLgRnBC8XLs8sI7yIua8
9/xZsV93v9vuP+CrFZvbeiuV2+hWKJLQzh63sMn2tGVdvWClkh8moiFMQnQgDkvf
vq53BPZI+e8UUk8Qupa8HXE8eA8/fk5SnybdDgE1+PMX7K/2Qp9a1t6teO4KloyA
uDHpv8S5UN/CL1birA1bhziyXFlGvor1dMnauQA0pf9/4fPAtqfMhjMAmHUt7oUs
1/OT+vUwBiGSmJCvN8BehahIsDVl9ADP9D+jINcjQ2fMBj1x9Xwk10KzLCnOsL//
lUcoBOg9TxIzB2/vKGCIftAcHgpX7JDxDZ6KccSSR4Mf6bFWiiE1Z24e6x1NMMOa
aBXOkxM/zaxqDd0g8N0UEvWmvcnPa7SmfFSLcMESaDPz4jtjSUz/faoirI2cWuVY
eEtREUTKj9D+sT5zyAO50K1dy0Xx/cXf73iCN1sjHfvXqfYUZ2e5qY3N2d8lb0Ea
lIC3L+kOkjGFl5A+nT9UiYHThztX0btJVDWQNCd7GVigjxy85MHmfbMOBSSSpkBh
me4YKN4GBeaIzM3ukkLuZwnL2xsYtbnCDB3VCrCmQ6C5+eKbTcnCjZ0kibcZWoca
CNRdIb8VN2o1HiFMcEgcwr3NmS8eD0UzGCXKbyP6YYSmbyQJ9Jwwpl6JbjS8GUDU
+pSyGGv1fKAa7CTJtNgPzxvYepP2I3HLlerwZuUS0IjawDuu8pbpgbrKsZb25veV
5wLCXhVUNhDGDEr8PZWRu7AvetKjgJKONn7g2mtm/ZtsUtlhxQJsGVVOmSe/Psr4
MTuFHR1+E5lwD+M0BNsILTY99Fob+tawiEvdefI7n32YQ0qEe8bsXDsjgQDqkpLG
vMDQ7DhK1mbv+Z+RZq29TKy5SsLQotN0xzKXINR035VE3uuqb+ioCn3x+11uBPLt
GRLPTzzM0FbzUmpTgbHJt648wkfSoAbU/Em/T7n5wq4Al3xM95gieDWSOTHt7g3A
waQOvL2VI2YahbcNd3+kLff3YMh1WLjiYk5W1dtjwFy2oUxuqOKdY4SuDoxJxvEw
AT4/vt36RleDBm3MI7YA9x55hBacf1tMvIa84WSS2oDu02NvKPyaaY0BsH9C82Qz
matpwLgIzY3Moix78I2xfjEy9EgilEijMuiq7GqoSDN4JPegG/ZE7BmeyH6BwV1c
RqALxStp9wZEYAAJRWnhmLnFRi25xZiO/MdyxiwFNOQQkyqWl9i+Q/EM9om+kq/K
+DTJbcSrnjZuX8vZsdFM4bdshPvjaFsR/G/EfNM/RQj4wZmJYuDjjahCYcGwksAc
HGtZWR4g2XRRp1DiCkrxXoX3AKpzVW85ik006LjTfzlrnupgTtVe4aW4/Bu/PqKQ
92pEqPLurBhrMUjIsOf4l+3vQ/81F/1R1k19ZlnUwVZD28DYfmAvsJ7Zkwnx6/MJ
8hPl2o//Ld8fLY0w8cmaZzd07q4mpSOCsaW3diHaTVXeW+hxomtyUmsh6mZgVjmP
33Tj2CvlOSY4vdWVvufjHjwjfTEsqlnuB39v80oKSnNqPsj4a83ADkhU/rbPB48o
fg6u+Ka94exhDCQemdAxi6UL2Ylc21jixaRFF6aYtmxC131oP8lx/zc5KMtBIv3V
TFJ6TVN/Z7VlchQqTMCOdv7EWPz3+kXZnhpuEPNADaBajPjzsIa7JHor+INSwzNl
Qhcr+OtWwC2udfM2otIA5N/rEcEIqgjoZjiabaIKUNUFPemNk89MztKYa3LpiTOX
M4ejfDDeSUTousA/vZQoRxxL1afkmsiIY5TwPeoV5VRkdIG9isxL8S5qT4cZzkE6
6qsrwEPUT79TALGa5EBK4c90THLg1RBGu/TNV3Vj6X99O8bXghXchb1bvZX278Wq
3nqvZHjGL9B/s4aotFHBN4HB6xAo9HM9MsGJ7n6n7JIetvv9MQ3yWB/pKyY6Ixr2
YtUNrDc67XxTOP3sMVQN9KpuoneT17zl2HtkTtmEr7AlcL4F/UYNq48JjkeyAMm2
feATWGgqK4spKFjYESng+blv0yrvil1zN6ETrNoSmrf6Xb1ng6Ys7T/j9uE9v2OR
mkv/VSu5nknEarEP24eOEIE7RT/xdMbxsIuV8tYcWCj2TyLhkq5q5hjZW8vvFjhr
uSyKRy8ASq5sELm1XK2Frw8EPF0c5LvzQ4Oe0tjRn7FbR+JeAeGpIHTUy25Qj0eF
yBH7Kk/tUdRH/9/is5QhjzvbP27QlM48Luj9bPs32/mlhfUEvK/p586x0R0k3DqF
pl8CMhhwiRzmqRlZG35VDRSLJgdXaPwNOL7hmIkNZLHrXaBR9HyBfzB/kAFVXQCZ
hefsQqnKMfZmCP/kGXCQ+C1pi40oHpr2bA36b/EaC+UnARTqchd/cse52/pQSeV+
2ePX1ST/Simae6aAKLSfa2RxPQ8bHevo0ueDUwjR7Fge0DMf9iSeJfLrrQWiiUeK
7+aQZL6bZuGSkhL1ycre8QkBfqcesIFP7JRbvAw4858WaCn+GKPDlVH/JzSgROqK
3wgKwjDjjrIFLdQlKyxz75KiG1OUOJKs04K3BYrwBsXQV6lQFr/htB3+jQ7Sap2e
dTCfI+kP678g8pPkc2utstVKPqJjMH6VEbc4vxRsCq9EYiPTxGk4hjaUHtWW1r6g
Fb8baH49ZYbYXeTshFpW5M+4/tTBbDWZedGRnesnN041vGVfpAhYiAVBkVKG8JvU
i6ywdNmyEL7737QSP2MIFEJwBOxGL/+iDU3K/GGNRlyrbJbN8uWfg+7mmcyOtWGE
v3LqrtNHc4nvQfoiRwjK2H5AO7GovMN7Rz6VAour8/KpHi/+ZwcRi3APbRx3bNMI
gUr4Bi9Ex3wRLGBgQzCOo+ReoIkVZXroHwx3+Rx7KFdLiacRRLvDfNbD+aEjpiok
RGWqtUN9S6tJ8CaiRh3E6ygaZ2NKzwJJaRKEPHXTzlLuQTrZA8tfxAV2aaJBiSyP
tTGtyn9GZNDeczDETo8e+ZkwcO/fn0VKUHmEjjPn79rnKvWJvQhuLf+qX/3KZUz1
Zxp+21b2sZT1w3bvrH3LU+TYPF51g1QuleQdqzJdhT8l6aFpZB6fTXDzpr6bYU9v
FCqM7NtICVV3u0zWt0wDfzOso1U4OJq6afksWMSZuyCsHXS1A5UFNKsHEv1TNhmr
s4X/X27sf6MY3Sk7ydrKXTHpPvCzz5pEkD2QIvIY18shrdqq3fPyhHNG+EVCdBn+
Py4dbjuIN84ETdHYrj6eWAV9mIct8RgUKQUi45oYjDjt+0gnxC0Be3BTJbSrT+mc
SXRBfP8qfnCB1LSEkDSfXEQJReI40f7GceHZkcKyMhkyd70pzqNr6nSsujzf+gJA
7/4WWqB2iInfj2pJvlY/LwsuCebofUTSWvuR+Zs0TzY9cH8nNQJUOgYOUUIBGmnj
bEZKXQxTDiDBq9TjLP4ajI+rSfP+UQHuVDd2kItplG9YGeEG4dYVlfLPbwkzXHNa
bJk/unLingWbYpchsxSZpMkZW1NYadTReyit7KfLdQjPoYWwh6twgg2iXwzz/rlb
fiqIADwEOrWaKKOVrFKgnl7zznnAzEKGs447g3iP3EYKDsImMTs8gf5jETi67CoH
7+qDNnaa3dWZ4m+0ZuLGOISensdZTbMQnHZz+S9RKfQ/YxfNDMTaiEMSaTB4L6ua
kjP2KaF2MOGvQpUcnqqKpR4VLE01S3gYpKgC4nv0jpJKcI8ImSxS2bQjqgtU0KbI
WkTXARBPLjGTqZ7ulyHrz5WgfeALaalgiqrKvtj0s+kr5IIjGpYxNRl0IPnz7B48
wTnYc+5kL5v5GK2ljYuAma/YNLmIDWfuH2tSH95AlmOiNdafPYVquq2bprIO+GoY
UXpIi2NPJRL+awAYUyrLzrS+DLJemWYwAr6zsqk31pZMbXp/VFKTLV2Z43UiLOMP
cqD1qI4yPP6hlIION3kRNluof+ybI1AxNreg227QpAm61z8lkwabYgbjvyBF2HSK
1KRHPjmLWzdPUymKgFtN8/q4MTuo8z2Wiv3L6Rt0GOMwdc7I+xkkAA5jO8GZvobp
LG2aQiXf84FD0c3a+5M8XeRJvkySWjf+Zk+sCOuQT5Wd3/daGbCX3CRRiHN3UaGl
K/w4hJDoCQr3OxTfXCkka/gxIf/61XAzkxanLS851YZrc4GdrCJLXFalK3oFjw7g
TZYwuJI63liMr0unNkxM9J4uS9w8KHsgXCOWhpiTh7LpcnDx+W6YCBxrXJzBtVBP
soR3A2kAb60TLX+8K2yTJTLM7a9G1Pr1w76uRAL8X4wPIilYg7vidys3g7vVKzjq
G5JzHVwCLN0RIYFeQXlfxcrD2XY0krJk4CV1V4rCE5fQ5Qzb/tC/sePtVcr5tvvd
S0yLdwJqCINnHNJ6H2mODlF3Ypw4Q+uRw1PNxNNrBusNI0LLRl4rZsmQBl8IxI7X
7faJmp3oQz6whuROSS2wK7wzvIZBQYwAGH9tPgaFypv/fdb61PbJkEgKFPyfHI4D
eT3ozkgLgV4KOTpil8tQ7Km+0mGjqNpX+cPDLkwY7C3S3Cs3724cIVlpxZra4NBH
+IVvfPaXpPaUdEsi6KmBjExZri60z5GkXrakztlEafghPJJ8Y//Te9Axt0ktF02P
Owsel1IZ91frmvSWUmI+8akBs/bTXMmKxHwe2mzB0mY9CSJcWSNYrH151XaTJxJ1
/nJP26uMBGJemG1NZTqq76kkZCgVRg2m6am6Epxb6/SEeNfOqcogNflpcku05/tf
5JT+0KWqms7AEVVwWKBkTJvp+mQ0M8+3u+kY7tNYRPpHbusW4S+vnvwYE5R7tY0k
uzsPCaZpAuYm9ss16dKbpg2UrZuSVDtdLOdwYnrd0IZUWnI8ju9T4YBh5CQhFGkW
lK47TUGlWp00E5FXS/KFMU0hfb4lmiAwMYS9+ZN/ZHM4ytEOabGmTIkaYIBNLlYc
fXM5oavzpAculJ/IJMIHI1esqVmgCkv1HEzE//sRwYTqD35oZ+Hbcmd0odi2IETX
jEW4U3tB0hkpGzzY4A7bW6Y1H4osbzVVorkqdArF/hbIN619pKxQWPtgbD40o7Th
ORcEq/leXscdhzn9wIUQl9NZ42w8MLLbQaxEOpdCSbjTJtOwviIhtDk3a+n7eyf4
xjaeYidxCW0y8zVulyhaD3BjBTk2NP2bsaDQSFW+dsybJW4bB04r8L2mGECiik/U
Tx4+zBObT2J/4R4A0s7V4tWota02t6te5SfhYU1UCF18XMCdCrWErqZulnLoNL/4
e9eqXVJ1n5nTyLpf/8ToS5/9S8Ajp5y4RExyqAdLQW4LZLYw9qcf7tjMb271dWiD
YWRvk3D2alp0DiB8agDArGQWjyYz5wcwSD2TGlMtdC5s8VzOMs7ULTm+J2HyoGY0
RNAz2Ipgj1gWIzhapZkJTdn0+7dwrjJUpCUxBDSlsMifgpY1CAcr7tTbjDkpLt6R
Xxq9KBksF+0NEHFP5RX3h743BMboYkevNsah5lKGrAE1zbo7pAhCoK9liCcKY7YN
B6t7X2VRJ/PgjRWKc34R36hxmIL4CgurEZkWlVmgPNX/NTlNrn8whNMZT+zLntBT
UkbhgSgHRujiFNZDdlPwnoDC6VVbznHxztbCUN1SK9VL/hi5vnSxvAKFVUCTM3WP
zRqNTBTnH3XaBhiXC+oWh6f8bQRyKcR+g062el4L7fnpPasApnCBgz2ICElIkURe
ixyprobKgMW6VUqQV3Kep42GgnxlWaX67oN+khKzCM3xdEYacYuoG/Ifwe8rx8ep
RJfKmqaNKDTmGcfFFCmpD0YAxidfIidplcDWcECQRABRSvcQ940Av4OClbCI82ek
HBN9RpaxtA16aXCmjdJlcotbxg7qJ5e5YVtxDCJ4B0w69bT7A6osNsn9NHosQ3Ly
GztpApfzS9DPcrFYkyfVagvF0x5zgkMKr5cviC0lRe6Axvl6K+EsRKQbflk0dAZC
75E0BvJDejhhPyywS4VUgqcUd8x20OQdARQpnNcU0owFKRYFhxmELXUVzZcBsaR9
YI2DIpUIC5tQbfUOtKrhwE+ZSbOjSLqGlCkQoXG5py2YCq7mlyt5BdvRvej+9phB
af8wGvo7Y312xIYBTRsfa2iZe/MmwJXYF2Igbx4bdC2UQe54uk0OjT7VAeBi16nx
kZ51mOjibxa3N56bOpmBIcmNAjR4AKLHiJdue/BDCm8BpdQK5BEZIMh8sQvDHWDX
/EQ/JigwOBJS7GR0bFX71gPtSpX7dk7DFfHv8E5rYBsemSbpuTUn+hREFDCEyHbV
jG9MXXnuKrljuPj2rQ1LTWCVfKAz6gk49+PYp//kbWZ9N1ny6e1iZiVSMTqJlB5n
cdfl1MC5jrO0kuonWPn8LHpWXMP0OKOhCdiv3fVw6wSKt3VK84apjz6ZIrjeTUSY
W/aACAYlImVXfybDSrO5rZAIupGRj2Zkp6xACMZB9sFWpRE3VF90P7DcwWpn7q49
R8stqhOXyR7tkAOLEB+8aE8jivSUebN8ZGL010l/VrvI/YSaPz+k8ICfLZ9Oxq12
d4Z+gXqB5j5P4tS4UN8oyVmKPJUL90p3v3ukIzgP1Dcpkfk4yYnuN/xPq4D1Hv/w
fey9kGTNlLNZimzew+FLy/DPNjdAL/qX0dmw29L3RET8ChdGcxbnE2WeFcotidW+
Rs76CBtgxxNf8MZHMZFdQuOGiomYEVcCTV6NdMxghLVU4iBmh6u/bk557h8c4/We
TD/5Agl2MF+mpIBzASZEBNOHZpqFbLzSx7OhwGNSs85bbwXfCEAz/Ffr/PBjC0Ih
iqD3CkU53lLkrYJymATyuS6rRx6haUv4FOhqqGRVSS2C9yACm5D3pcM+KCANGVal
XMFvNA5zVcRJ8f80q79w6vu1KOkxKLH9//jNRfcb2/xnjy4fVfbdbaPEIXykkXaP
HSQKfw1jb0jE4cWA+cxLgvqGvR96OjboXOiJIQbNN5hQGqajINAqYS6KqpShFG44
SDtFEjodhOYHXUopdXGbDGjcZKm+XMg2W7t3JBG+B9WwJ/chg6FnZroijv0/m0cV
cHiG7eJbsKHdkUdQBjQxcEtkE8UazztEz+2WnBKVwNy+jX/o3J0J9cHqzrtjRXmM
imSOBBnzg4jPGqhcHiVaUgNIYZeWTe0fBkg1+kTA34AFL821JIU6GR5MbmGvq/0l
kGbGmD1XeCUdD57+AKHhW9wrqF++hcG5VoCNdANds8X/6NRIzguU6eunlRIM5kPD
MGMCevHrsqYOcx13QNKRXtYyDO+XJ/HsaZ3zIB+i8j4Z+nwpgE+g1pXCHzQPdfgf
B9uV+EuI5G4VO3on4gz4Vc5em394/xh84F8qpulYP5N+bK9fO07SA+uHEmSx1+N6
atbKUoN+pj2yzH/tnxl1xts0EBikMYoalaCob9hnamvJmR8SoDmHY7AKh/9yABZo
+F6or+1LPOHgmQYaTBekRhSwQDqJRpZi9+691rJh81QE2wGxmjdsVIWUI7135+rB
h45HCZygo84a95RB7L7LPLQh0p18faQt8Bktm44Kitn12kj6qP+NknEK6JBiyJbJ
hHWOCrSGsOt7ZF0YxeAIaXLrCKbBs95YoczrYlhy/LuEMfMdmsLUX7HG5IZEeEs3
ak6U9/tq2uVlAQJ0eoGVtTIK1xHvhx5d5ZRjmNaIipq2W6XXm5Zcmc0maQ6tALqj
7w/wkniQzTP+yIhKLNbMKS1nakpCu7FAJgBRz24mkB9woCTBRWw56Yc5t+ia2BpR
2PCsvfRUXYIcC2Yf94cdZc47jtfVLNBtZxdBlRxnGpd4myT0Gp5gfCU28uNMxrKa
o98T4vHBmM0Ht5Z32AUy78U30CSxE/iFg4aFRQ6sqtO5FG22SaezoB0FtgDIHyS2
oEPx+MwS3vSV+k90GaqiwG3eb6zYr000d9zxSiDW+FLS7sSwkQEuM+YYSDxNHg6x
iASqB4M1SehDeN2kboKzvN9G38JXcaqIshBa7XPhZiqPcPPuhpvaRUxtXCg+Wrqr
oIy4oWFbgeTkBu6kLbgutooOBPGYStPrk2GyPtW3FmeRrIgm4LOmw4B825nD2Hrc
fPhQEa9J2mb3Jm5zyBCaGWT8R+YPyKf5+J2LLq+LLM46n+Od49AY2XlO8p2IyeTh
cySnZ7vviS+weuZL+moF0ZfM4pP2TjMAzV8Irp+nBoildQjFWwmSWMffDYbhl6Jo
lGaX/BRLRQev53bku4mcKK8xKYgkc0HqmPa0ybFR7Zginb0A6CsGxnWI6YXu9pgg
p8y96jyVWbRyQfIYWAvX443eHdegzvWJCF8wJBDlHO7KYKiVHp4U5SsTwGDMjdAB
qUUTMuN/149ZQaOsnYZ+49SSdcndh3QBNzsT/BvwlRgsn5OSSK098U107gPws968
c8QtrwA23rkekXnFE3LJZhjxr7+nXHEyEiTwTcYFWh6zRbKUXq5vXdK5pDP28yQ0
MqmtTw24+0xn6KVr55471WK58SxXk1+a711TNbUWOYuKRN4kurzBDSkytK4KCakB
Ui7BUeyRXhaprNOoAnCWxvzVO9+sPo60U4a0+eKRboX2hWMm72FTn/GMydARcIZ3
hgRhq0avqvzuczCyIxUyjdBGavmAUo9cciSACn7kaYU23L4+oN/Fxl0my4lyWOOC
kHM4fPPoxESoxiMiEfha3iPLRIQfNgbjZBXyntaAy5u8lgnSryRgTKd/1izwJej+
uCYbX72ulE7ZKTt2KBpuKsAnnrwCTr3Xm+B5aCumu1Sr1Hdn4RFm5GGFu8Zh2NAp
PbkWJju2jTav51rNd4bv2x8ZawifeBI0Ymhi4lS2cGyjqtLNZgtJhbxg448e2R8m
LgBYh/A18k8uDDBkWhQllH/BzbgJBxKyTDxJt9ulV1HiRHqx7T8M2VjE188+vcoS
DlAPpXjAdnJLLW7e0B/lf4DmYwRt5uKh8n0qe/7XHBu5i2TO69lno//1+Jw2gBm3
M1Clz8VknQ2yr+iSB92xA6cAaPygrExsqQRn4xRnhU0b7tbB4qXrfM9hb8Yk4K2q
Dz2Gh+Qj6CFyPwDBUZvHRmVisg1/rgLT+vHYyl8QUKNfZeVYcp/5Sh2bGIG5Xe5K
wBVlegPAkKm/ESrkaP6mfiJt3y+7/EXd4BGP8RvdlNQByEc9bWpkOqWV9qLtjAOK
x76rLDm3XuRW9uyPkjlmeBXdvGZfiCkHgfGJX7V8zFcHPL2k5oSv9zJs4cjcREyv
ULgjvB7IMIjFfnzEWMpgg5dfFSSAszD3lIvOCp+9FPIHxQ1yeJfMpwLlSLvYNof8
EOhMEAqMyOy1gYdAT+CleK6sTjXAhiwyhLP3vZHzauLsBI7LNy8ICX8M2p9UF14l
zP9k6O7sfm5xVdlyJlkHCGGFM3pdi1oUf/NmwWhu5BjjvaBVS3BGvvHfZfgQjOMc
ZxvV+ajBm7rB2QyjxoJAaKq3c5/VaWVvyTcOxQ8DRbKcp62VKzwSu0U+fzrH2O7N
2yFohqvIb4lhKQ0GumdlVN/s5GBmCGyou8OFgdJyEAYgTCDQXXnmgvnq51WVD0AV
bKpKojjX9ZSgZax9366D76p/t/2OWrCxeXRotrOsRiafaRqXX0IwbthAhCTw/nrf
8USEIPg4yUdSgCuZUdIcs6W8lmC4jwzd28og9dTiFIuWk8uGHJ9qfxYep8Xjp/r+
mbcIBnWeMCGlmOEUi7crZA1jDVKoRpO1lI5lRMEAv1N8ocF/wWPPGs39PRpVRAVT
ZCevs/eq3D/U16kzAtxucHX9IVsM/OQNVStuBemyjfGdnuBNOADt3QAC+lcrBVfS
551zZLxwGFgZv7TlNijZWjfJGqygf4RuJ8j+9fLYW/vA/arhO75tiyqmy2DKVV3/
IFr906BagFesumR7fILfQWpJoRKzZQiCYJYusuOwGcq3tmqT9mmcjSUfVNeStg5A
kKabN8xU8Qvm3FPS/Tn1+Jx8oeTgKoWHP4VAYLWCmSvJEaeL+t7P5P6xzPQRnbCb
9qjRERXhiS/23onmSFdOGn8we6s8g63ioltigF2IxxakGN7Qw44hdbq+YxJ0XsGW
YL8xmPAh28X+hAE04RfMJMXU8jZ8t6x4YPXRjGYHmmAxvvJq34V9jpz79KnPghLG
335ngMPWf2okE5+vMd18QLr5VFyMnVbqBs1kDjjsugikeklKdNXwFykOQL1gs2lf
XewIE3P9ZDuISmb94CE4ktr6RUi+WM9bt/wN04KFbc9yJzcpB79Zv3sl4zQpdgau
U1oAT7+F4k8gj2BzjxJ/zUgq0s8UC4qCBV+sfMcDz9ksmCz3CVf7u4HupOwPLjv4
a9ficBaW7YmGPALnw7eQeHdVO+9JhZRXRbnshFodGdDUpgylSjZlwQGo06lyU1vR
g/BbWQXQiwrofEerkKj3SDqN3C+96xEYVXSWiGy9FKFPJjtEH8oIAbAE8O5QiN8R
q2GzeyAm396GluBCMme68vHjoEwjNMKWhK9fIwplKgbxgAoLylnA8xBQzLYUczrw
P2sBZwrnJa5OsDqAqfsFcADil4jatt37IWxplN6GV/riiZFm7ACRic/WnNbnM55b
pQrxZvzMsvCcd8PpKIAvcw5ORqL2o28Y3fBhYlEAi8zra2DDGG9eE3+zDrSffif6
+e2IlrjYi7puWNkT9mXhv/snIHXqFTmxVGwaVTGnJbeQHPBNqO4EfCZTUe8hUXPN
LPGpPuv8fJNtocdPEaeaScHu4/bewzp8DAp6oHeOzlIsRUc49jAmgwEPq6q3WB/4
fxZTYsxNIXbXj3TcHCQHAxvReAZv2EjVrPr/hOCccmhccz50VNcxXHc8Em7MI6oD
AW6jAuD2yftDN5AqQ2iJqIgnsfqN8IoK7gnch2X1RPCUOCiXgkbP68G4JXuTD1tf
qTu/3By/e2TgMeg27HTuN1YQ5f/zmbmiJndx4PWym2Pmy/85y0Tv/5UrpppcG5XI
PxRWUK6nHg0yJrqs0k57zlWq5yfdtChibkIjNQgU0aevo6+RSwfENMEWkkVmsgst
ldul4cT99YwglCkh88gAFaSboVdNGZVBqEZXfX4tE7tgLBv5/sUI7CpyooU1g518
8cw0lcJb61i1lCOKELRpA0TWwU/ecbX5vEnUQ0X0pAnAkmRYuLm46r7QLnzq3uUS
BNJv1CeqPa6kSsPrnXAuAqXt+LtLGeDWTcczGsqqGkiYxaOFghG3mzWNat5yyDtZ
BB4y/mZwI+iZWY2J/Te4X8hAEAV3NI+W0O6uF8bBy5rbBFtdrFKkL3BI87Ja+DPa
e0fvoPtl1Wbc5qCyY16T1UDAxK6hQcYRz0tVqkfJUhHIqc4ovY3+MhWZQpe8z7G+
yBVrgG/ABqXukcXwfeVloZj1rAl/Q0pZtlptTbRVb8pUpbkHUPKegm+sfJToJnnJ
ABf/7ytXwjFWp+nUjNWmpRvIsHt8f4RyyOG5jLCbbZEyrheg1lP/Q5IVMitaJAZL
EkWuvr/OVf6QUnU1KAR41w75u00QELPgCXiG4qaz8D2J5M9f8pkvIeB3OjUj7vO0
/X/4LcmL+tyeoe45ER1ieYShU7RbaqnVcdcRol9QKj/1GZehJLoqbQmBACWsHw6O
4cBMgXj2GkMb/eDoS64UN/E9bhfMCIsGi3tm3QfFFZLsu/MLS8DlzIe/AXkcx68e
lqZ6Tm5dHpKe8A83nWhp/ZqhuODxUdHbm9iC3/EyM6XVX19YzATdp97+CPLKjvRv
qQ8/4KtIOax1fiN7+1zNRHIH4DBJGD1nejZvqRe03A3/szTo9HwOe68MUwFZ7i2r
dbGrpipBLMipJ26esue+wqjLM48VCReScPuhTDIJCpST1vWBPjbXGhzBdC3GUuBD
piQZUq5fojLJ70JZt9HOxfUtx6N2nvyRho6t2Clt1qqzF8yzCnP88aqn0FTpwrxJ
KjDBOTFBWHISgCWoArdz7G8ssfl6OXOhTESwNd3UQxqxvdbTSoF3QMHyDKsNhZfD
E01/HCwGSPFPJEhNRR/A4QHboUV2V3PFsY2aFcrg+oJxdzAU0eRJXTtCYrXRxUI+
1gNqOzvTbcAbSZYNOpPXb4693Xzkaw3uknHOsKGQcCUYM/ZsyQMtKDEac000zzCg
TP5o8b95disxqY2AKaEBL0e6SNM7rUU8fvkSCaWc8M20iyIjTL5v/WCx0zpMmq4d
UpmuYvm22wy1jPjA8htWJeIpDO8j6Slxwc4KB/7fDe8FBbRszubmybWx4clmlZlT
HJSsKu7VYR+JQbDkS+wOrf/BWsCCxKDSKj6y0DIuJjDfDWEFoL+mjdQoSwwRCK4d
r/3PhOU/pGs+NURjjL66QODdj/1mUcSffkwTDIrUPOYW5nJSzW/vO+wGI9IrYa6U
GfNnVVgVyjDIr+nAM3fv6D1N8lRmL8IA9tDkGNCqpTEt1DTTZ/pfudUNrOLVmsqJ
codS5V87cloCnFjl0nUxFMVc8hW8syMEOw5xzU7u66jZILZxc48vGfDssNExpjDl
JsQUHrmoTvMOaDlK4yEY4F0du8KttQ+nqln8vmcsUMxK/f0NRvqhYqSXEb2oRUl+
UqkN7SRCmq+h3J6cs5L28Lxgsp5Ud7NaJYTXE+E8Pb+IHwpeUlYZ47+gWrQfuiqS
zktRDgtIO7s9EVaO+w7dGCQkEvPsPZkDNObvivRTwvPLhvpQ+TOcLlx3HfTHkMbZ
cyWu+QOcqi1pDXDJzgMA2S+03Vkw1nwRmpIA7KxpkkHU9TkZDrcA4kVxr5LHqS9U
YrC1QwD8rhfVVEYa22gfyUsorL/yz1363uQI4TuiFC8+3HtlGsOzXpFpfyyEbYeJ
ch097PWkVXDzewBFcENSH3p1Tq7DUZByzjKVflXxjiZUbMY6+HwJlhrkp5iWjtXR
bu74fq1xuVzSuMD8ZCSSb+dahBCWBI1sahJi2BdPEqXceDB6ryHH6O+Ol5fUcdaH
HwEZlpT1GS9Hu4QzfA0GW7efPjgx9Ao86UYY8pftNyNLcydAgZEa5NLvTuhnIO7G
wtfrFfB9Z0pu/1bDtGkvVejNfJ64W0SX5NmcTbilljgk7/28pdYgqR5+b7KbTWRe
CJHykS0VCxxnPiy8tnyJdzqvcU6gdOWpZUkqxCZvT44OPmhDjp3KObPoaUTZaOEP
9lr5zW4znRZGkAs+27PE9SauDidd7KwJakPA9D0ZyV/UFNk/pZndtYdAY5QwNqNw
lquMVTtXGoFfVvofszoC9wbDq7yhp+tlrIts4vJErSvp0ywfiGIA1Bjo2DfmFAyo
n6iOTaQ9uZuk6quxFASEErf7cRVPR1O8VnYP0lBltQqTPO+p12P5zfrgozu2It+4
Yi/QUWmtiRlz42JrxgVsqA3JC9A3UV9Wh+IYexjquDPRyLpOwHCVnhK/gMBzWazc
AQcO11BAX+9rhIxF75ujJTv3Tz1LUYGHE81d1gTS9jnfUrb9Pj3ZCRUuU2Y16v4j
WxcrtzZ13e7LMUyw7xSe/o2quQRWiZ+yJO9LnB0msYQ5E4IocU4HfqLGcSGSMzFF
HTc5H7uKNWQK8DfB3K0G8QdaAT7nLJ3m/NYmVen7gsC6xOezv65T5IqLP5deARjp
TVWm3Rr5aSsuV2Hmk4SsVjUx+B8BjrlWv31JctUA1ideMZj64uEJBPBZTry56+6n
UhHVJn4VxmKtN6E0h5TSBRh/v/uG+GlLEmgg0X3ZoecMw/BjMnjbbOUfhQ6FauH6
grudXg2m4d3XuQBkXMp3yF27qINQL1ewG1Q4wxFHOtqZPcstheZnhQXxNFlqFrET
bl22N26cAhW5GFD18U6tjRKbfo3rlhKXYbM1+3w86EWUqoE+5nhXMt9mSC4jnzPd
Ge28cJb1Hcd3Eh6uFOQx904wUwsHia5UuA/AUELrODy/eFlm2H6E8Jraw+9CsMsf
cJ9SdnI21/n8+MwfgTJHYP7bqONG/CMBEvAzMwo6GS1/NA6849XfxfaLM2Bzq4ba
L1g3eRzSYVt17lRY3nBU5AAUJZZJeIZlrYeCgW0nMTJThqWYlt4s3Ldj6LHzF7i/
f3ertWG+t3riG8VVf1X8JGmgW5OOQkGcPDhoCEfraCJmUjsZsM+sT1KHdAVdPwN+
Jh3+ytHkqFg/JGCVH/noDKStvO2uP2o62cOlJBr9LduqQ/1uGqbjWskj1cYrLlSr
dU6WYoi1DFcOVWGeMNaAys/ZJwc+zykbjNMuc5zigDbOO+djDc9oo4rFA2RhgjCd
A5mkW4MMyJLCzt5C5TftcurVuD/Qf5ka6Qgoms/kHfHAEczfmo0SwxzpaaON/ESH
q7AOsiy4KsUy8BODWa0BsgP1aj3rOd+WDOUu1Q9zhVHp9B57RfYqr9pZBCBQhIvE
U71UfXLXYY/Xgw+wRXplBnOxeTWBOQqtVXquUkRurJ5Ago/VJpDCKFVgS21hRGCd
UHcIBGavlZfM4hGl6PXGA0miKaUiFpY3kCMyS+i5jDiHEy7ehrd1vjabIFVFYtk6
TT2cP85dWKtFlIGUE2QU/3b5E2q2C21Hs7SqgKh/r0vZ7I4mpHKrXW8s9tDVI3PE
fUfDHma8V19dm9kDSc/1I6RMS0kaP0+c65HX7HmGxqQ6OWgIrGa8yi10eslk5qGj
L0VFeZeTPveXC40e20OtYTB/mDbi1UiFaHUu/p3xzG+Etx/b5pOusnVp6EIWTrV0
wk3VFrN8dkphI6OkC8mMOpDcJI6HKe4MuBL2jZXiqqRdWPcQixjJEc/ofN4Ura3L
RfJwpkoiOxEaatvofxyOrTPksFg1WH+bTjF5dh/9XMXv43I0sEKQ9ogqLZj2kdHu
taRRsX8/LvP0IVj0L0pbgDPNucs+OMKLtXgxmPAzldwPuHFiUzIJE6ElFA1ldyRQ
ji+D3rjI7SWWUMT9FXpYSfCQggWB3B+2psxoNEZ4/p6W7lZbwhFBbGZbJz7h23sb
QHa0rKXmhYjnWuRhZLvdpxsdUm1XSu9DcwCW0LudZz97XT9lGuUeKBayU2fpjuvK
/me+eH+MH9b+P5lJdEmE5GBtDX5//A+hazjkSko25gXRJLNCVW7wEEuuhQHo91WY
UMyfJS4CNLctZDrLcqGb+epf0j6iecVAesWWwBKaOQOEgAfWwBBDFbHQOqIEsOyN
3qCDfYl5NaLBLgxvrmy4cnbMVk6UMqHEOevZj9NAjd4d+CHaZgcY+tOcWMZpL2FY
g9+9vY6WpFHGp94t7pZg9mQb2qyrGojsEdml8hY7IQ5pOQ2B1XqxYEazL7EqcFGz
BC33vH5aAgBQOXWK3dE020dd5OsJXXMkTLtv5gpq9JG39NjIspOkzpejanVA9Flv
xHtZWH0CuBdfrcwXz97w//PMZyXfvYJQ785ZJ4p+c0yMF0uE/xclq7t6KrN1X4Xa
GeaIoddPiE7W4jiUSgEBUlpPDVaANSarkynTosHH1shbyW4Kn2mIOFIwp2czY1Y9
phq5WnobCylN4sTbIBdWeh2ZQk54R0gyiMhAIy/cPO9tgj2x6k3wsx7JQ9yQ1kwk
AZ+xmF9n+w5nGsODY1D1E8E/qS6EdyOebaqsZRjVluzA5F6CJN6ygUUg0rI2U7nv
d6lufkR8KHYtvNTYBTnEfcjYNvvzYqlSTlXte2YfBkolkgIoPEK8WP+9RqP+YOeU
KY8pUubNwcafbpxtRoHVCWmENkfCnEGZy9fv0ajp5rTDeokIg4YV2MZdTHnYwvEv
T4kgtrpFHVY0am9FzxjMZfd7rjaorfBatR3X4sqUaIWE+I8y4rnMV+6iPsoY4du8
IWYltUzbgDmo9jqWcqDYimWTjlp0tLw4J1bZd8Qq+kcuPnsOHwUHNFmbj6eE3web
QWxCo4AfQ0yAd4ZOHxFqWZIRHQKRtDHuNEZljXXJOsl4sVkOSj8U+wrgRb2guhn4
BJQW8Xi5WkyrTngYTMRRlZOGMCrdx/my/fyMC5IdCaiPC4FpgeolsXUJwTqPKzgr
tQIC4XJjnBYnHFFLwpmmA/8N367uNhwk7AatOzzS8Mdphpzb89h4EKfr3oX+DVQ7
gQvpuyEqZD3Q/RmbBUI5vrUL6tBu2sEo6y95fw54loUyaEtCNa7cXiXLaqDz3hMH
FU0jqYoV2AFpW3drGs4fXaYPKLr5T2qbMsKa7mW2WTaCX7tfOYB9x29qzYW8AKpP
Tmpw/5rZNNXmQLdsJeUIPrCrElKUco4ly8x6Es5As84PqXbfiNEmOMpgcN8fdmTn
7+/dzoUiSv522mf72WnKPvKu3JIva8P2Ecr4ct7Sv01uiK6g10pZw4t8tsf9KEuq
XQpr29pPtBv/0SLFKsvX96EAV3vhWgQTUS5IMf92p0DugtROjSJlyphydsSd6yJv
vt5htc5d+WRWan9L6Trg04VWnJ2PJxtHXGfFJCdDM2UAGPV4mZY5uyn2c9S/xJW7
IpPFDdDQC2D2TXmqBbz7FbqDj0/kQGff1EQ6zcYvf8vHY77cj1hfkufp1XnfUXEb
3+JiaG1Tki2iA1hPyp+9xaJH7BxLOLb2z6nO9okX9u0F1HSLicL6bfrcieB6ydA4
KYtodwMHIOesrUfx0rI8xF4XocjNXRLnN7msS3BuXW/73VM27HJQyl/TWq9u+plR
sOSj11kQXlYvKnAf4wBME8MkeO6xns0UovUAM5whoomnDVOwftc7Y/uvs7etW7R2
7ViddYomWAHI24Y7MgmseJk7t0bQ7P6LHw2Wub7FkrYcNXGPyfbH2vFzzXvkFpL7
2wsLrU8ujwEHBEEXBQDkKQrXQ0W0IHMB5Khyitd+loFUYwz5/GVUmShNWm2vl8Uv
LDKuwQKH6sXQrHog2vsif9OyLXYj3xnwtzwPYs6VLO5AJedoJku6cqsAH3pbPF/t
mMekTvNCzUpPppDLwri8FJm2YyzK18wQI/EvVS4BODbjdR8y4etqxE5CjDxmTdFC
YrDh3tkpcoCDL6umUMdl4VWVzaU3EpTmGPfmEfO8i1QUaLsshnr0yHYJPjHokIb7
MKHvh6TbXxSqlbi6zpZaoo0qUPy4fTNastrKWIUZQ9A2FPTpwrMv8ENdhRmV2Vzv
94DjCRNb4N32+Di9jwOeg2FyithuB009q28iRu1NKwtXJhZC60biMRAilUseH4ck
G37LN2JyNz92pgmzHSS3v1meOvxTobSxOZ3TZwXa7Og5lgkR078jE1KNGOHqpBsc
VafFNPxcPrRIJY/Aok2675LJGB1lT1pmFSXvfGn9vyRyTlL2yQrlAqmBR6DyaUrM
B1rjzqA/RO8p7B4aGFq/aMrIgd3BXhiPc/cFgL65XLT/tNy3smyOXU7YqOW9HUUn
eI7i7NaNpGk429AR+AekwrapWuye4JlWzcvvsI2qEHcDTfSFJLsBPGhfM+Fz/gCD
mnM22mHgtSIn+f5ElIX+IVraTel/PYyX5VJFWDWg/jC2sOl2QbpVriGqwsnW2cPn
yem50rQSShSBMTZRUacOoCp0No4OMHS+qAOuIXZPEjPPuAemRi0guDqoOwhvQSE5
nPYJTCJB04bNlcZIY4CpwDX2GRdEqpxAorvukxC0ffvS3eY6zu3ZP2OEq2VxkjNb
MLGNukblwgvqba95y1wtpk7n1hqKMnCGFeTEcnsUOii6T29wKG+b5E4MX5pD7urC
XW/VIhUlhXZAL6ImKV6PFTb2jaFlPVazxiRxd43z/nqKCut+Z2Hh18t8M+TyMIcK
1mSldf3w5jGY8IU6+TVSHclkb+WM3Zigo7/AjvuXBKsOn7AhKRYATbUqVpxyexxd
h8iXzsbhx/cmVB//3pRWNk/Ujf/OMJNkSDX6X58nOu3a9imslOJjpOf75TJSjQq/
nzpz6akrJbm168rR1gayWu/SE20/GQjgQ+lqzLpo5AruttG7GFsiomf36nzFP93/
Ze9R3qwOEQw4SK8bzPa3j6RIR+4tHRuHUrOk+IHF1WY8JHNOsAEN/58DQl/ckbbf
SMd24//P4T4lch0poUcAwp2WsVdEMXjvirHKlMPE/uZ/483xSZ6BVO/cSqkbVUfV
qHPlb6uQVVL2dRRVTSZovlkEX4JObcS1bG52T4brdapBMB18ip9QX4JtBbA0qGXz
pGyYrK97q18f5Ddy0IKHfHpPfqaBgdZCyeSAjDBGB2s7uaaNpzlXjVjTe9bjTK4x
dVUnwgU2B2zgFqmVAy/PlbZx1cCg579COEf2gY8MDBubPozjH1zfAyVxoOWxB49R
rXg/8Z1T6l0bpLTf7NIZbY+C28FrPjpfxUuWdGrLWplM+sz4jJWBaSjKIpKlTZj8
6U47wtnKVjD/i1WY/li5LK5Nh3pzkexE+RD1n0lLqoKsyNNeMyKXofOd+gCTXr3/
R7LyisIe/eJ9d3C2OfWvmQEohaQZ5Ogcv3GB/5eGMqTQq4ph/0QJybrWTX/hMe8O
UyACC9fm4HrQEn4BTUdsYb+Pes5Vkq4lIsHJi2+jYLqv4I5fCyqdz+ZPibSceBV6
Dp+++g5qkmfyPUhAQCBhTL67/+I39WXDCu569ef4byz5/nRbUeZFPZiJHas9b0Gl
o2eorKVv4iKqAMWmPA4Nog+qCdxfodBPEmNRyaB/n97q2XfV3bRZcTIiqR2vCuGd
x3WTvzh7EPtVxGXexkOrc1bBxg8vkRmBCYqfpymhqlw/WbyUEH2Wh+uiu8qUPCze
i+c08yAQNw/k16GFZckZwxznTpVFgkrs3SIKPfG5EvpworMkldX/ySJ6zh5aoxig
U9lZeWFCsKgsyEaGmoSo4xEEduA0va1pTDxnFFBKo2MLRogChbSTLJjEOLJYsKow
X6QcnEWAAwFC0RJretlj9B0nF7mi73PL88R7fhSyhDSvJVPm/PWmRvqpzk8ikWbA
zcku0e8nc71Pqs9JC9U5rDB50Zt7+zAdcu7socdEoSZqipMR6UkrR3nkvKrLFFxq
MJp0GhzN6inod5LxZMsxevdI6BmPvktBnN6wGfgXMscXqNHln7zH4B5a7VdtfhMz
7/gZcvMFtxeWyEjAA+XG7Ea4pVXbziXAtMiTV5xoIEiNLOMgPCexK40xAEDMY7wY
VOWurqHSplcnAOUgHq8U0jiBPtNETjuj+aH9PAXCi4IRR260fdg0G5wE7aQ0IiTq
XhwtucMUo5w/Kk5NFkA1Jf0k+1EBc3StW+2+skTaCbFOa7p10eASIT7lwHmEQNkX
88p9kFiSQ0z11u/CgVrUy4qD2yFOMg4W0UEQdILtHLGXPy3AiEHxxL/0hylJMf3S
ZfkEB5W6nSm8nVjyCaemCsxOPmWfvkOreU15VjbAcDiCZFGW4IC86IYy2FkTvmW7
46Xcy9e4m7YAqx054PuknzGwd0nhrGcAmGtl4jlyMjnGqMaasdzONNh/nEt3/ZRq
7ANtyUqH7tntQPI0+gzZwaak3K1u5lbxNxDGsYwry93vUlG0FHNTeNvVqrTFaJEP
UlPvBG+fBMxFk5RzNBGNQ6e6TA0HnGlf2d+lXsxcQgAYjjYQhlhmPIqdi9VX86uG
SgBRYiWNb5EG/6x0C4UOh9qx6n1vNqf9yu9blvyNl5I1Kph3uI7XTwY57C+Q3Or8
URqvU1wbsr1tYezLW+Zi2W3heFSXRhPJ+gauSfbph6vN+Jyq1VViYUw4jCjT/Cao
uBepED8szxl6RGCuo4G2cbRMi0Ue4+zp2c/WPjvPKJ+tPQZZjb0C5Y2FRxiusEFq
ixp9/Xjf4XSofSnpcTS6gnjGk+ybGUf8jE8qgz26LlgaL33fV9YwQV45Zu1V3aIs
aZn4TtylGdOJpy73HP7DxEcmfG1CTmUWleLYgGdkLEPsOXDkTV8II6IaLGibnZE+
+5kD+Srz41Hzybbw28AMNIpeA/AxBrRXShxJpICWh7StqCRyMkTcIGcyEHNwBMsI
eVHAVZuPM3B5xrobrH+9tS3PX1c6jmOk8ybuWaLsZioPvNG+FX9cQe02v4Yfi6/Y
acT0fF3TKrcKUrlH7ZgaNYWH4t9krSCm6CChO0+Jx7aDD9pSzJqM0clv5jdyAS6M
RO8oaPMakBqu2aDbDodkX7NP4QqyvRT8i77EnCRwLfqp0Kvsr8srSRfIZutokgvl
Sapq9WVwVV1sRm4Sf1i+cMDCANQBLw0qI795iTKcUoNCDTFz2m7Ntw32PTsRCpGe
Nd8OzQrFhr6Pq5oUhnUZ0ZW0bTONOtkSsU7jV62m2h0GWEzpOJRKQB8i5dMGOSQV
30Xi7AuRlFqnoBtd1ESQgfSs+TpXCofgaVntYYHFUdE5KrAPIc0eBK0Gthns3TsC
APaMv4dFMvI/2hWzEQjc2YJRbuY3/ZfeT02uuaCUyrpUlKnqkl8vfAtQC/Ddqvc5
Aiy/kBQTdPwskxQ+i6tcJRkY9lP+deTOcd9shoCDW1G+smcjlhmNcvd+YKhLtYhl
4VroA6w6UpB7O/OXaxkcbVEl4cIQiHVV8cKwRsf4dXdvPjW/pMmzMf7emqo43pR2
3PFo9xnIC4kkSDc2x6rPBHuEBUqZ5I7DTzjEUjKJOSFwTWzq5MQPfvJFBhOXtIgr
RQ4k9/ecWbVZ6OWW3dxM04erVH+nOtStjBWbSPPvq5j6j5dgjPO5P1lQvZt/UqYs
ivhVQrTtbce20tlVexgd6U/WURNjBXWfNssql1KIJjUZtQKCqgdKPtzmpWJecGCP
+0Wr7OHdrRW4VFGOovJZTc8FdiGqcjwuPCbKlVS7jgSPTuAgIhnPwaOhrNPhx7cb
wqwQKi9MVjfnJKw2/eUgkjgEtYZrDa9FU19RneIDTFZ0Bk0SrUfF8aRZok24UKgs
NYKA4ppqwQ+MjyMIRmX2gO0rgxE79rYxwIJMrKBTH60Bx3daHfvqcYt5QaOMBGRG
ZHkwS1DLe9EuPl/ZSd+Dmnia2xK42j8IEhiJs8okLl5b28ABu+lzQ+Xqup9B+QLZ
EIQhbzck3hFVhMqSmyKvcdkQmcpDj8ZYXhQgUEyKXBGb5AQ0+8XQ3oGwpFmdL1ao
aBP8qXuDAcvzJWr8MoipRKsX4ULr70IvIz3L8XCvCL/jutar4Ln6+S95370MK0rj
McJsB/6IzUqKxuX1rUCWe9f95eagSA+clGdJee4bHdGff8IhGleYdy/8T1cCH/7Y
6rOs5F0ui7k/XukrDtvamdRkgCYCAmEalarjgZsmfRr4mXQDXR2BcNUfYHqKGOhU
wWDPk3bCTpHGBKnCPFYoN3O7xPpQEZDx3PmK+NHFlK1T6KYlPtSEH/hZRGS6toG1
QfSbrLu5/ZcCINF+lnY+C3QSIKKjVKd2g4iL8o/l2mhcVUstqn71pkTOoDuVEBZQ
Kj2yldgb+8HxszsL+PfcSS0wLsFHpNJCRpydViOzp6t+qVIxj1TZT6bbPdbPRI/3
ZbpejKWNwIg2KGMAn1oezGafBqJWHCTAyg7/aw/a9oPSz8A+xGZJrJKU1exmj3Hp
4BvW3Cqquan301GyYr8R6/nXYYGAtT6eE6vUmQ7IJ4bIMm5BBRRGNV6KTv5+RowP
PxMPjy/1vS45bpMMAKiGygsubnWiX2Kjb3PeDkz0ydqSNhPzIEsywgCTy8+/eKud
ukoJBO4VPZxlVRgVWMqw7GQFtgNpscE1pZFuT708m1xM74Abxrpk9hjgH9kiuEXG
WFvMJ35E6uC+e4svSE3OwtKcXakL99iSk+kQIlZuqqjBwHOevL4ffezo03jgVYWF
+dCkHmKlhvf4TmfNnt2cKInG3lQ/sjBExEhzbyeHWdBtCPg4tt5P3T9nnOSCUBmV
h356KVLnA3nBdhDWKxtBJViLNnuOI27i5gNdPotJi8GSVrbDgq/TlXPAiU9Z/7/L
Qmvfa+sCd8QZpXby+n3BM9+iTV8tVJHJnvJaRjAPra+Ssqq2bz9BqX/fCy8WKR9r
OWDLReDRQrS3d2fuHM228mjN+tgZ5DuoG4X/VFr1FCP0NXodyhmtOTG7PN3F3NrL
pGbiG4dV7SPx8yGBaNxq89olkm/u4BeclWJufz77s57FsJxjAi3LhGDT3chdm8IV
aBkxA/2bAfYDhTRvEZnLDVng5w7gMdEbwtyIuOuMr0aI7VFvWuvTuVSjlqzAJLx+
Twvy1YH03ZGwhm/1H0C6Usc9r5hPqyHlG6wMo7l/q13oUIJKrJ6+MLdn2m3vvZBv
GGpalMBBfOYkHombv5g/bXyq6qjXov5gixy+Enr3D5MpnDte4rOr3dkXWdQo4NYp
sYD0tashrA/TUD7IcQsdi6uKf2sOOs9yL159kCsCD36LJHMh+TTbOskYtEN/x9h7
2qfDbKPXWwwgUULT3FZ9OB6aWmOjJTeilZ8mJqSkx3L5IXDXHsggahJWGkW1gVP6
yAtoTlqTUD6xPnuAZFPuT90XJghlZ2LRwk0trS6enFP7yqDK2E7JOKCxjj6oqL08
Brd+k/ECY2ednD4NQHiK6PT0uP5yYCLWGXR5VQs7Ht2/dH4iD5hjgf7tQYXth5nx
SIWxHuTzZ9xVCm79ENwDIy1iOEF8AQfV0h+hTMHCAsYZTHeI9Nug6nlgUHUSoSB5
Eyj4IrvzOs/uDEI9xG1tkpbPSdb1BwfTWYySYJmUXwXoIk6bTDprjtomBSR7UJGW
MyT8TCXiRmwcuwZI7IC6I7+Bdh3K5YqlawLW1Z/k1SUQCJUdO3jZYx2fn58IGYt0
xbmSeXJE0M6haM1tEwyx4YwUDcFfoR2zLz8Hh79jy5ZdCdyzU8WLo6wPFP3hZu2c
mZkmHB1/Law8Ftqkhl8K3Yk2Mh89ZZhKFOv11STX5LZVAP2sZbOCleDe407gL/8J
ErODN4+Vwag1kwRKlftHGlCYDdOC0p1ayqoooCx7SFO6VL4mwOhO7/OpIDvnW7Oa
+oL4rfYvvWo9uyrLbHR+DtpqUz91PoF1Xe2bZfmSH3pW60yxCX281VMEkY71Mu5u
FA4rhJljlPo1fvIjxQfPOPC2L9hwv2XAFLLJK2Yf//pioik1yuYKlke+ApvjSiRw
+6Bbv+A0LnLvI/zkGA/mrUSsBKUYHssf3eKlqOibv92+ZOG8q6oSgnpYRdtD5rOu
7I8k4EcoCZRwsgb75Rj2fk1HOIlPcE8zf5CF0dR2xcQSXPHbYjSg9U7UZXsU8ksC
VizldnKOmNv0pSCmMVRzIqYKSbQ7KSGAh6ZyhgDOrBNKr9Tq4GV11yDkX1E0IPuA
PiNG4pgdMBntI08dDtTR6afQuXOfVJvIcmEixsEopNNXosQUBFOIt1wZ/t8nT7lo
BoQCHM3OfWjY8QVwCwu8MkVzEJkSfnSpYabqIV6V0fKSzMpap97mKrXJY1myMzqG
RY6tYLHf0MebyL3dRtUH3WfFrffbppSwNpf5YHDEMOw0IgQKtNDhSKfYOC++DYly
UTL3DjhyWbRSPYPVRTddVdGp4lTw/3GKwx9T9T4jde2W3FUnqBFVVGbykcbrMyvO
LyjU6SFs1Jx8QQps92Q0QfxFB+BYiBbHk+7U+IQdKNPzhoU7XRyC5CGqBlSAJKYk
nRQdFBeELSS9/0oNYbX2NS1F+CQUITQLGKV6lYPavJf1Bytl2HQwwETJ/A5wOg4w
r9c4YLphGYX0edq59MuDA79ERHwRIsz2/MsYVOzU8U34TqLf3tXB8wdMqJmCYJxf
FwWc1SfxLbTmTXa34wXl7sjhP8+vYietl/EkLExiKoNE20Q4tHN2xeiDYqPG920E
tgQedyi9MAVLbCjT8xvAlymCkBt7vTQTE2Mhc0Aj87nOUcW0C28Io8G/sHKr+gyn
SH4fb8Yxp2RX+97B2tfiw4Z//zRzu4exQaGsNbs25o3KGZroTeWq5KcIvlozOPtX
IeYuT+eLy8vn58fmkjbMXxzI1OElSzVI7+kj0Gr29yUv6MJA4s1/t+FFMIqqA+CN
id2ZBDheiDmK41K9bzRT9Tg7xkKsUzVu4IpNQOer7odnkYjy9RSWvmE/01ekDnoa
hSvrJeRdLHSqHcEA7CHCknD8h29iyFEtZpAwrnXwDQCQqOwIyW4lWXzcsnHgmM19
D9p/ja6u0O7koMS+CoQ0WHvCa+Vy47a7CYGiYrqdhsxhjZuNSoYREzGw6EaievNQ
zEiCtaPsnDFx3k3U2mMHNjCU6zz4gyviK09f1QRjvsUiK/f2R3hZq6o+9zdxqTio
KSIk1R86iyZsX2eQpnVngaKsxSrVbkon6tcXG8yLe7yqvgoPZUe2W15PGvZzUYo8
T1WSixEgVpcvhv89eee9yVAcy4E2VvoongIcDlJslM8smChsMu9vJwYeHQNmsS/+
Ymcw0R9qUzM+cTyb2cwUGnt/0zEGvvj3SxOGHQgn/U6mrShLrEPzIEFoli31NNAt
/8XilNaSWF0OMfnJZZWoNNzz66UbCKCjBjfFcufnXo850IATADf5+gnDrB1ePYz1
7JwYkuaYp4SKJsxoDhjH2+u6KLb88A94pmBMEC5Z6n//hyWIDTRi2uY18aUlCnTo
40oheTZMtQHo39eeABncwPmrT99J+kWewz0RB+1RBdSz6S83bqf3ZF64FzU4n1lu
NBGynivRRxvG/MRcgvwIp4KrDmaGSa+IlBBHeG9d7LzlGX/O0+rmStG9u7HNb+6V
RRG929Ff8Kzpn4lvFXP1YbUrVD6uV0SaZmLGRxebzYI0rNt5HW73Jm89J5ahuxSz
qNrvxKlDCkJpIDKvHxLj9XPu/rUWMEaJsFAeKPtXfKUX0BrNwJUARYs1XzxLPxHI
Nh0NL5b6RCTZpX/kY13LuzBQZ54Prv6yEV8Gi/EhMwNnEyQBdqhB2NX+5te4rSe/
qJ9MuNuGmVdL+TwpXmvWl//deo3weJfcIt6nOm6noxLMolfXQ2PYAsyaFCA1Jr7N
OGqrNTMYI79wy8JUPFCwcMOoe0bNKcSX1L5YWYdrCgy4PAQYnlnil/BDVNfcqXR8
RYaMqlmHgRmzH2LC77rXiLld6SoauZfjrK0LyClSnmxAjUASV1DSffGK3tJlnJpU
eUtzeBotAnEvv+y3Lt235h1OfIaUVUj7kl58T+KlD7Q/8+hwIPT3rjEaw7RPYgBg
FIOERGhZQif3Kt0MrWXNpTXYCUqaZkGfyxfg1qC5gPPMd7oeWLgWYdlF2pK2sXlU
bagEhwfGAfQ2x+m9DHkDKrwjSk9EGsYLqPzFwoXJPFaUAABGYVUoLTXqYpb26+/+
GCb0SV7ORLtLm4uEceNEkcYLifoKlwALfQf2oWctLRENxq7+rjCl8ppwGioMaSYw
JrVCMU0sieWcHEGOSZPHxccrv03RqlV5VMLvTABdHCnnNrN5RGF7VNbNfslGzrtu
eTSJ6r/DWuh2Hst7+H9BCmdFKZTng9Pmdv7M9cwZ+JdfdEPK3Evm7HViFi2nxOCq
XeXHkZOvpkvkLwTTXu2567/+rFyvKV8f7l3jRxtPrzsIYyhxKJ8m0iN3CQGVu/xD
sTyJ8bCS9+pd+189nuzQ5+XqB9kiuJ/zmeI+Fhoe4UmvMj/aVtRPZbhCGvcYRoTF
5vZ+0E6V2V4TN94fu+oTLvyIUBw3rajy37cyvfKU1v8CDOPgpZ+aCpcdaS5z1RiO
UMKvCf2kG/QgdqKiB0larRSwgW+rOY73TaDHCUJQDpnw+LvnfnV7DrB3ha2wkmL/
ky0fkGTVYGvwJS3mbx9EJLkg+aRwfGn5F7aC9XniihsYPOZEZYgPSADm8zEDNBIJ
z+GxwV8Av/EareAynqyHbl+mBmEVIilsX4nUww0V6PXHmiyJwd56tLvcnXfCsM8E
JWBRA160IORsXPthei2U9G4aswRhVA/lfYjB4fXRSwqDmysZt0bVICCFp9NrCTXh
jYC2bd1ZxGr3aX8pC4rDjSe2Ssh/yQNDtEhu4ebisKmTiIv7zJTFXq8kS/Z+Uold
tL8u/j4mnxw9KhSyDVK1qIoxEg0devMlV6kGr17jbi6KF5kL/VTFK4oKc0AuPp/V
ZiIsEgPkTcLDKJHRCVkgcNmjCknGKedmL+4r3N5YwBTUDhf7Qmbb9EB6u7pWz0yc
CtRQ4zu52AfWQQUdfFwFtqQeYmWSz40nGlDD7TFKFHi/lVKJ3+hOIqvrseutJE/S
emPrQ+xSq5u3pdnt0LoQPduuczA6RQa0ZvByJ4a/xjW0QGnJQqIJOo5cnBtQshW5
U0e6FM1CCzg2sNu52a6w14O08v6BJaoBhyq9d3/SzHORQncifsc4EnQEgctJ63Ni
cxenJQuaweAKSB7PmyOuGExlyOygd7HG/PLqKMBnS81/cFlomy3Jg7eFMMwlXHvZ
ER4RI6fQPzTAQOucZobU3P4uXrqa6o8R3W0lVDijZIcPEgjF8iJzt4viGRwOZVmM
oN5iSEs7kLZ7Lg7R99RHHq+AKqcAiSJ64Ptb3lfO6tUYALzo++HMuDVnO4YEUFIC
R6wjKXVG7M/PaU2oNoac9oulmYvX6E2ZoLcD4q+v8Kd5lML8prZ/GZkqUiWE4u/Q
m2vilBg1MzoP/8MfLKvVMFRFROFDzgWk74l2UmFO7S1749vycUXuCcxaKf/chSKK
ntxC9zPQSwgZYg+UTNxkGxuUvcvVzYT8a/LmgxZJfFxkKGTiTmb3b10Qv3nGlPNX
WapPyYBesZkvj3YkNWW4Hg62hGOc4nZlcMpf7+3S2N/7l06olh0amYFKs3uMUYAP
YNlx2MmJm9g4Qho2Ws9BChJxzbIo6P1uy9JxqIldVYphgofaJDC67lr1GOyqlwXu
4sNf52QMy7LLLiF5xIJSrhyj+hdVgHYJxPwXAKqR3xpsPehkBSHojuuwO66rNUeq
IY1l5PqP7rmEfeRZi1Etp0K4GQpVYtic6zzxoo1+0XnvnGjM51h3Il5Kge/MW2QY
kk/YmTEVJNZgxNIw51nZbpRtJK0HQR99w9XcAz2889TAxMeph7WATWQNJYwSyzZL
A2fTFhj5wWkUUGojy3lwloOiLpxkvZpOC//ZFceAFRMA02UFOSNZuTa9GdZnYXsl
C4yaC1bt9SewoE3qcvPKgyriidOD/bXTFiEDRBe83OhnZJ8Zfidb4nJ/UIArf878
pFLZabQleQvhhjzBwm/2FUjwzdVf1feClqYRe+zdXb1LNkOrhBT5wMKLLRNohXDZ
FqyCYoUKtJK7Ya+simrbNmFH3v7d3u83G/eIfYmf9phsczQrMwPqUpV8ZtpvRskT
UXbkIDSiv3/rwb2+xQuWj3Wz+DSis5q+QNLFBG9zTxbHUmDA1UZs0T3QqGxnfz/l
YViN8he/51iGW0g5A0YQBq/urMbEkwig3vaxR9WLMehULwobSk29B7YDIIqm05NZ
IL5HFMqkh1wnLtpH7ZPViNy0C0k1XSWkq6lGtkFrszoyl+pPgN5f0JrlSbdFeTdj
qtzcXb3Ex90dEORCPxqSJnenT4sY6Hd2/jpKUrWrszltMXIYz35eWD1bWGqT0TG0
+7SRPxoSpD0skU0+XQbvCIlAT/ihhNnZg/2mRbBWTt4ZLSGJg2XnzAliTaY4F94B
7I2GGmnrwl8mt59RVvJwgxOIKa9lSOBFcRe8fPqr+cwOB3IS3sYIUYzirLlu3+/I
Mhq0gMEH79qimrDrVi58qlf2WYCnXbA3jEHGooTM/vGNYw+cqdr8WTV6QmQabHRz
SHfeA8SWPdpXmM7CD1OcO8DRsIoXzqKmiyMF9RwDNNbKPEKXWu1iG7vT0f5gZtkj
gyZYWpqTDNPYzvXzoukDPlMsvw47GC0saRS3WkKnOvINZm1Sg3i78fl08R14WtB3
t5jTVY1Oo69H+etEFTHBVvX0g/zR6TUUTHt4+eHlSnH4fDfTG21RlCI6JdoGLHDp
ylhpWIho374h7qj6rIDQxDpX/y6s2BeQ3vLrV+0gz7RmN9/5bLw4yIhpBGNfDSAy
1Y1nSO+VF+gb0DlgIOe81hy6TqorxniUE5mNJcyTQmr91/JB32FtN8NROr1YeuPU
cn8qAq8xxf+PwN4ANwdV7CFrpfvuqWdNLQevL9dwwQUrwoVPlIYytrEi3ycc8Ufv
3sz1p3FcmWtSxBc0Fj5dxrTfyffC3sueCoLQhieidOwTAWJ2IQpnRdSRQg9YDbYH
ZSOhy9C90uwFzasn5aGVs2PppL2G9Uv1GhFnnCPvQnyiQ8chUj8GzWqnADPqnvID
a7u37TmOjuGy4iYLymVqgcPmWzwiqqAZBy1AHF0im0o5Q0WgYH94WM3mUYx4Dvvu
hQAgoaDUHynI4hdP3ARke5hYH8KKaApG14//BLg5jDtCWr4Lb/WDZXdOXuaikCKV
JOHr3/pPR8+XcxOQB+9PqYmpMz4IxqfA0L0xuLDJ7wSaxD4M1ODSAWRtuBH9v8I+
Lhcjr+REqwCv3dSbL+bfIB8kEIRkCYgFwqTh+GE+OT/aToCMr9TTtdd3h5kHPf53
/ChS/i7GFQfaNzu98pjPObpUBWz/90JxjKhjM0tt26DyNrjVVJog7MRSiwfZBTDg
Fgb+euwdO7GVsc/xnUSANxo32QQh5dfYuLRCdhD6jBYu1BIp+VonPANGIa9/fJNm
HC94wsZqU0jo6gWkCVyw/LKdR7dQ/1X1iv5Y+V6PGXCE/FKWEiGS5GHV/KWw3pjk
C+Lnz1/x3A5R5wBtu70JB2KFjtZ7HV4RjaKQvQT6416ixVoy9iCPIE8PfoJ3zL62
jFsIjOhqhYjQr0cfSAXaBzdTLkoUMDk0TqPklriPd6F3hjTcbjTisn2040WIsq1B
nTGVGtRXJHiaaAaw/qqVvj2f88aukqvdLw3TbsAWbOdkDfjUhQVoEy5xiiSMvEeR
mNNfQY/ULYOa0B+iMK1bkkr7zhXCnOg686MS3wja+pgc2Dkj+HUOX2Kz2vjT5JE5
7rHu96A3z6XGo6k+3xJG8ZUE4fOVE/UDFF1V49fdUgvIJjUikHoTMwilprj7pKaG
C+bd9AWXMA4APm5VpkG6opDeXSXc9JOPQxMQkzxlpQFvBGEcZkwFiF6utRXMfFN6
KLkZwzWUF15OOKHe3Mw7f7ZBvoGe52dd4ipi2eQWZAT4oi3cQWwdE6tADYLgPUJy
UTRfxGneoZ7Py8bWNiJFhzqBJroAIaNlrT2Z4mPp9fxTOixe4CWvB/NvupKA8se5
qI5OVMWp07TQnFofQiDJcQeJfC+4lgG39LmtB9XAXqNFON9JwzJ9gKC3zrfTabq2
dajVJRu8zreNgcrhzDv9AwvaxL/U5yV0e0C0JcuaBCRv8++Q6MYIID8EVGK4SfRG
Drn3tpzTKwY/CBPHCiSjvco0wlxhZT1BhKO7sDBHyAn5jgww0F96WPdmnTHrRiC+
3kS2bogKSlFldy4cv7ImpI84aLy6Wvlbjb9GPm5h1pSjQXrPh7QgkFNEbalMDpwm
GT4Cwn3Pv2g03hQ+f09UVKejU7k5DQGDozAvXcz39PWHJUIkFtWuQw1yuwOhd1x0
dsljlm+U34/WWk0IhVPjCkBC5hhaQoxq7aB2Vr5Kr9cuaBiPOZqin4zRrhOWGBNi
H8HNTqSeJXZSFiXZAYQg5yMauTbAj5toYVyL1PJXtouzcx8TG+WQtxzzFmKh9EG7
g6UWRy8ohfMq4jf0/mEd1keOQ2JWI77pgnwwrkL4+C6KxVLX7cDb87v9zVj8CBkq
PssUva28txsKzymor2nL35nxb3KLTU0kx1Ax4aRwLJg3xpTmv4fYXzXDV1+3Bv0v
43/hD/TsI53v2NxBxyuqL9yBMqasXiN1R1gN0bbLIjIxL/tSPANMEQ1f9pMXQvNf
rC7mYE5sSoJV0KGBjh5do6v0jooI+If7DaxqExCFMKvybW0IHcRMhrnNKg3Ucu10
m09RCjcaDlomGSzgRpaSZ7MVoW3KSWO70HZCjk+UfkdZpv/Ea8zrPNlN/oGJvQo+
n3R3WwA1huHDonEV45n6Blp2I+Lp5gPqgVEvPhDFZuiy56kAmFozWK1eNpXaNnDw
PKsi8+BSg3Bct0hG0SE2gOMYyxvgTBO2JyR1naDUZqTClnrQ607hhShmXYCqxRFa
Iq+6MKzUTEcAg/y7/61DlzE4Cd6ay/ej93g9gBxbzHMkN0AE6Ejnfdr/mvPDkR5V
xkyzWmfopb5Vnqqx5SKMqBJqM/HDFsqyHYzA3AUlCHyX5hCyA5pe/QeyDH8r+3Cf
mCKlOgdLiDCsCMJrwA0mKfRM3Opqaj4zKlKE0BkWotN0ikzhxjA99UBoYMtGaTYd
T4+vNoiSPsVz2Z4AC6LnTbynXmqLgGxTL0Ba5A8SKOHH7U5BT0+okf8ZR47PArBA
kdubMoklvGIsEjoURpVgmAvzFsyyddZ/mlCP1iGxse97CbgeeZIKUaIDRp1WRS2D
ot6dpPD9+xqY+XMvtazvwAOz7LSUMcyctZBfN7NdJ6LVsOQKJVbwMxMOpUIBaC8m
aj8qDsRmI12amBN+ZOV6WXIHuwWQHq0iTahCRtUEXcQID8QKGHhmNqijlLh2Vc4S
Q/BXS8BMXNTeg4T9fGWHaIeFguYsSKKhnHqmE2wNNJlqJogHlfp3cxXwA4oZ+RVJ
5WuTodbdAgru5RKIACwuSDyCNTJcQ0kgbRWbNnIFJK72DycoJ7aNA3+htQEnSsUb
A1Q9UGLAJi+Tj1nm9bNnX3nZLtDzVXnPvpKajjALoUKw+BgcJzTA5C+qIApBZHRo
bA1piodkDG+ECm2FIWdCPKjTi9h0NHBUUHMjljc0bzgyaoi3QM+fEsqqvBbCvDPd
iXCuT8rSUyzD6DbNGW9Guce4z9ZTbrpHNwes7UJIBkzl0YCU1COGumAlmt4VYNL+
1g1v9pQaIkOEgTijnz053Zb7F/KPmDa+UH4rDUpj0WMA1XFf+SoZMzMjTnOA3//6
YPV0sX4qCnquvH+CUvsCXBlVc64MdJ+pwx4L+aJ6OUx0bF2HWoCKt+7ULZDNKmjc
MnTIoGHjuOyPlSEXt8UonxED7m6jelt7fBb1D82yB1InjrxTz3VE+/aVx8XmrpZl
VnMm35ey4r2fZkT8GgijN2sVA1s0C+tO7XEdpsXoXP3F57NiEjSzdkpTCjqsNaDE
LN2hkawyZZcVdQ2Pj4w9YBwy8eVomqbjX+Gt8YdOJRsqAErjMK5KN6apH2pQwyGt
6tBoopG6VaZ8/gkQbm55QGPSsXjVSBszQfThquu0e19QYXwzHjcNUJ8xjcRP4PEr
r68s/prs3ZWJ3jKdcqiOzRXoGW0gwPDMFEL1H+/BmBRrOpMewp0lfZEiirKdBqmW
Q4ltXWzOsbWuPxfpWEnEgCZm+fOzkC8KPj0C3iAC9ALFky69Xu17Hyyq5sl9y7QI
F7eTXYneYZ5dCMghONH4WPw7LWOxRfo16VJApRDBBQNyaX4aiLT0VhRlTEndYmwA
ABmlNyn3C4S4AqAUspC5Yt17c58wSrdpeJ9ck/mBfZ4UYXKQwsUktmGFUEGW4cMp
ZXeFuO93iB6Azig2sOKzdUmG1X5im1NAeFqG4sDBrhWMutU6OdVRVua1buVe+/YF
WqKFDTxkj+8cVtOEecTCNWvZnNriuHLhzn/3crI1jXPriDchRt6+H3xVoLg/Ks+r
ve3yyTBLfWRPLesmT0JNfYMXoOASzP0P/nC+dRsaaAxR3zsXhwD4BexjqlcbGqKj
77G9iTE9X1VeO0T53atxleHPtWTX11jQvn/gn5otiRx5eXu2WZx0BcRHXbDTRvbS
2JZ+VqJ5hbONaUqk+Ov9NAagHs54tvz2QObMGt2jxla1OaxwQ8msJuB1WiwGiHBR
zn0hoidPmm75IU7EPWiVkHWOh20M2uh66yzSNcDc1TYAXaAspQKo9QQbYRUFNlRT
dkbN29KGLnz08iPHS1LNJ/pgfKrCC4IK3nysxxmYQGZrjtYIreQHjFdhBNaY6EKh
FxDN6NAHQoyBkPe6b56yg/9VTC+Z+q0yQcc1Zm22w+TqjlvLRoccr0WF2WLbKxO5
dzWJ0SEtzXiX+U24V+SF1uG6kudkJEfWn4BdZLPzTLZpfHR3p1kvYsFVgSdP9AzK
ZWdGfa60PvsCZ2eiMUmpAnKGLS8oMfhCQCMQLvGaWoKnowGzIoIrEuhfz+aNzcxj
soZB0DVnmRF8si+NGeu8CYxJ7swZ1bLYtVfnv1jvbgjHjqEMnVpwcVeKFOSU3Bio
oqXcVaQbZMXKELanbnPL3R/Ir717WXlDa81RpOTa5S5PZoQ+w6dbJ+lmrB1sRoXG
8cSjLcPrpu7nl7d7Bu74oTd+JnJONjdLH2yuLASf9Bb97EvEjPxbptw+ZmOnfuTz
qK7U5ncj1sZX6Z9hV8FmThqdXuFuUyj+1oabOXZM9IgQVl3CtPwqX2/inaHysGTA
wIpZ9ntMhcyIPCt1QflqsJcP/YKqRPJfmUowsjNWGlHiakFtsLPfiMr66kjOiHoP
HCsEd2QJoKXWzYRsl/mGvAVE5xtLcbJC0Pc/iIBz6zbxw0WT94Tvnm7D9huS9Mh4
OgzG0MYl67xUPkVUuj00hyY8mv//v35sYqPoQ/YDJQSDemgOP0F65tTkkGmjh9WC
QGgR8agLHQanwu28ArnkueEsVCenHSsXFKa8o+bR+iOaCEA9MJv4MWobJe39sSRV
v+8ztxXkRwQcjr2+rXXJKh1zDBYbYRV8tslw7t+H0tyqyXIotScU3tjw3Vkhm8k+
1/hFI4N5DBhgE4rv+KJfHSKXygIQn7guZkcrXqkPdyvlDp2dIXJxjs1KSWepYmw0
y1/1CDbqcbEnodBQTqTny4ks11XKlwIoNHD2a8N23dHtUKSLyjEN/Uw9+rR2dKNb
SaQbvHfxt4DUmnoKXnkuOLSvQTrgTZ8cuhngvS5YZJKvfPWxGwQGmbAmxjf8bThs
yCQc21nfpCc+4ZzIFiS8nTLY5tOqvbe5QtNwhv83xJgS9wN1sq0Nneefem/CVp6R
IjiM2WySrHN7UHlklsGFmaiCEekt81wo9iB180VAASnxjCgkvc/ofCX3JPViRwOs
ZI17ufCKiZHhNGDOSrp2qYWFP9YNjf/cj0NGvWyH+QX/Rw5RGKB8JxoBTSLMeUrN
qbDtPf38gsM9pOHCLKhkiufMv80grr9dFrORkBuWIlt1L+WmiB5IoKsH/no+Ug5W
byCsABY1pVW3uKL4n4+yH39rYopP5E6KHUYOzHc5g6R3uKobN9Bfa1xQo3ga/sHM
u/2erfPS2FyrP91q0fY0WpjhqrILf4kq4fCzVepuWD/ROXNlQHEuNx7ASFG1zsIG
UWrdeTkymocgWAM85UNJxHvOSyEBmnSAm6XkiTjWkM3+64UoPD/yeGsAy+C+4NBw
kqzIbdHf5/6v7UyAUX+lE6aIUjXDiEGlf1/jexJkabMAQx951FutUBiMwf1T2EZo
Q1uC70HERqw9gnxE1tl8i87f1v6Q++OYbPMAjSsJzrW3TBLEo0wXtTX+EFai7xch
oF2cdgFq1nDerHAfPNSXJ19J8q95bORjqVkN1FVWqKk9pYjs3CQCqcOt8Ahb878L
llbHrauk238O3wGbnZyWoq12jCMl9Ah2qbNQsw4rlGiRbtm3m04GMJyWf0bkyYol
ecXuTkIbDBugg9DziOSGUV2cUnzY25+MHW1ekD1P1j9Z6rTJjBY9wLn/6RK9mHfR
de75SoBMI6xshDTNB9GYN+Gs3rXEJvZ7zZKKvpiqfB04xsFWI319MNjemRbAxHb/
3mMgMFt4P+FIGpIbV2ARF4JwKEv+MSu9fXwQ1nZkydZq4tvfYWMZZbbUmiVEKkk/
QJM/o2xspqiS8nMn0g5Uob7nFTicAEWxmST3PQ6MRKlB+hLG5ZBeLL3HyI2pFh4b
WPst0z3+TpCGWnq/Bjf5Omu3N/m8YZNekxS5vuRzUBWR+ZvOIUCYlDkKZknxPfXX
G6mvyiFt+I5QHgLtP5SwoGn1NqI1VtxchgRYhxLrHxgx1ADW60ggOLYDEhD/9nQh
1E6k0/VYJD2fEuxnChLy9HiVqCuIBGGuBNJNomqqeZMK49hO+WsfQRaD7tOFOZ/r
M0pJQ6G3S1lsFuAN7hhkuMec+Wsqj3rG/TNlCGlpJvzOBjhm6LEAo5C6m1oRWhBh
cCDR26tStC/6TAKU+s7lrqSTZ/lIeogqRe6cBHDvdV3sR2ssnjDGSntay+cHRdXk
M9VXzWk01KBkMDqSMMSiQIV6z9p+8crStJOAN0qxFN8pcHO04TGOlgo2s/eFd+k8
GZF5vMOWjnH+fRsZcEyNMWJ9gADYZvqLB6GPgcHlJJnkLTTj2c3IFpgyMdagEJzQ
r3SKlGXfKtr07KsM1Tlo5jqoLDkMPPax4V72Qdm/d9Hb3y4ZLhU+mq6IcUm7yGzs
gRWw+2HLBjkbF7NdpkuvPS8uqKt5+YZ4FSrBMWu7UtmwShAeL6Uv1NFNBNAmbFVX
WTtpXWiD7abx+xTGYNUgP/kkN7wzn6h0GNuMHWBmCrDnnvHW6jX19nNoVOMDO1QA
UaYZC/4Nw+aH332haLeqExesOS0Sd4lwgPRImdYpSztzaFoMtclcaabj67lqcss4
k+cHes/T7SBHo+A9RorHxdr1i8yGN8RfUcYdwH4354aSohbEIb5wtEXCv18Xdxww
0gSE7fMtnMHOMoJgx1/5RtDJrbex6aB5Y8+dRp3+ZufUyqvZdUZYk8fWv9Ocd8rQ
Mna45fV33IJL7WqBD6rNmyVGotM0tiU52TYIQ6MT7BGc5tMLbOHAPRvmlZv6tf9F
K1NbG8mJG6O9Ccs0/GiIxQEcEaR20Ut7P2BYu1UMYUd+MiMM3i7Bvo0mLXZ5C2TK
aKRIRZvttYBOBC+CXufReZ/UniqTEd1c6UqXnVNjZLtVXXlTV89YmTGPm2GqFpt7
YjaSRxtjnnHAOIpI397sKTM9DcZgLrrAMeAhXcZTLRWuTOIEOfMYLjT3LgDuD4/4
82USgCnpt4eF+Zid4W8zoDkSOGL//kQFeiPxiymS/SrGmPVJAzlcVgDnbKrrwHGj
cE4HZDQHhlc2tSZ00DL2dDW3gOkMgT/ZMY/T2sHNgvTDv2i0jizfczqW5kT4McCU
6D9r4aAdqjNVWd0r0XzPXkbHtNF2LlLGTQqd4+c9uEBiTjChEH16aW+60JhcKMqw
rSLSKUYJaJQpnI+YEc8lTJ1WKm4YPfJRY4Ls4Mb6T6821oJ/U8OINYOvdV41KSWR
C4H1TbPW5nRMIebGk90P8xwedha5UfCHjMIaY5eDf1+R1RSp6tQ9Sb1y+mOacwz3
+qTNE1VbCR7C3lhN8Hb5KD2hlGh7ZHoF2aMvYK+825P5u9Ox7KOKCItIYPl4dT1Z
F0f6gCm9wM9qD/PvqKuXa+UdzHFH+KxyCesOGPcgJhCEeXxKiFk/Zr4z3QnyZacH
UJMmnCKOzx1lE9FMzLLbP7uGx2p1hkBG060iNrPZAP3P7GOy6XVXO9DrWh/G2GDe
nP6LWbKciP3Wk32Aq7RoKq6oHxesb9hdNyHyxcWT8aGjiwxJjxYik4nNPiZtRfIE
CQf1/ggVW5FkSeXQfrbTSkETMawUH5tbvsRquIpAdPQnr0JQ+GmNvaMGwVfeyDjA
XhF2YfqlX2HbV11HurE+gwN8eTIUxm1x4nFP/lniweiwCBogsAWuEUtUyPcSp5oQ
Pq33oSh7v6RdiWQo6rnarBzpsCrLNw14vk1twqY/R6gT5eX7+B7zOb0arEv2q6Qn
7IqOqb/AUnEeLAVqAT6edYjB/tPgh953A/LlLRqQ7o0pyvgfaFlgDbrzc+vRcBfK
yxEVoF8iy3uzxsHRcgBh6B6lxnj6GJJD3Qd3PvxZyjxiREhiZd0PUzvQbbXLnX81
Ml3IHLJeqN2IQdX/rI+QBU7zHwtR2XGnH4zjqA4UfRcJsG8vufQ4fdrA6qRdhTw8
epJ4fi+PralTq5CL1xo5O3qZ/6DCvUY2QxqIyEVfD7HC+cQpLdVjPXPeXyDDGa5B
w2pEmACxy4mAiZGDu0OHFVmy63lMBAHeOFdD+z4MoVLzTNW+yIqm/QsLSmh0PMt2
WYuPKbCioSMPgpTDN3jeCh5tmtRvbJkziN/kN/m/785ZVZ/UhJpku7pGByAuCx8s
I9Vq/l+uV0YgA9K4J8QXJJa5fzxRkvk/AhCFCcHyN98Sl9cHGgReE1tbvtAnSJOC
Gny0k1m14IimOfXmhzBP7Sdl3JmoUCSLXXrvRBL1qpFB6HiirmJHp/+Npw1roD93
1E8mQyssWlpwu97ytd5RFrSfaNdrNmUZiafY52T+YTu4zv071I8IFMTcGA2VnbkF
xOc4xShpIfT4gM8vmta0wfNUVHqXGxsMbaFvuD4LTDejBbyVNt9qBdINIDRPqoKe
pHNfbwpHH0Iml7KdcJHIx4Pr2MI4posF2Jxr7XsZdvU9kyeR2uroWO/UNUMCNe1Y
8rx4iFCm1CnazmfYgkBstNYu+c2W02fET1RtT25yU07uKJpyhOjPOYMKzvq3KxgI
zAu3y3dfJtxzIQK1C1qnpBOIbmxQH7r50wI9r5092X19Fx1/MaBegYIV6SAYKkAE
25xcMRHV7a9PomrX45w+V+NwGZByw9NcbERiLoBctTVLM/RAWlNDg6He2agfCZB5
s8sb4XjW3L/6x69nugfMFF9C4rD6VxuKyKLFxFKyW4aKZCLtAY819jZ9fXCa0bdR
z4x+PUgwoStRW1bx4+fkNnSj/eWLiEKD8F/YJ7l2GsZOV2vDezi83/K9lQtzZKaW
JR2lfXAuiReXD4p+ahf0R4j+WFW7hh1uTqEjm3rZ4RuYTvzpqMQMyJBK2x7SyQD8
W9eywwk6U9pcIF0c72BX+gh8vF3cDeC9Z/pAn9HSD4YP8aAT4IZVoHdlbGxQek09
IdYZjidnYEf0vfitwN+4m0NQVRIRrBDmN+yJ/TV2H/2z2J0VhaA5xCMOZsnDjzly
ejL4T5trrdO77HZJmBInxUKK2fJmjOdIaR2FaCyh1XntzWkCCHZ580cRAmfkuNai
knLFeO2WecEXYDGFeHbm/Vc0axRtVeZ9WRayUOhTCBbfHSH4TinIPX9FfrLpuO8T
1W73AKYhtkEX8Oa6kVANEz6pGmyP7/BznW9+XpW+aw2jdzJ7zprP2Yy2VWYVBqZl
Bjfdynr6JnZhQgTNZpb/XI5jSeo5RqMtuJNRHf3sA8k4PASkepO45nJ6eWoeWaVj
rldIwazmwnltb6sx5PqVoEgPRcvQ3+Nc6KFZuvXOEQGaVGMy6Dgf946jQYzqipBU
XPM8Em1cZkGAPZBpXJEY0YRr31PftUhXzPlqXlnbQN8pwbNo6fXk/wzBfqIaXViP
+h7TUyIosbfNLfDNvMHLxaflSbGlnkBdBBzMMnNl9zfuHNA8n2mVEw4QKSKXs8ib
TuCOTpTJdxK9u+ouD1EMX66DXpoKLzD44N1PQkn2s87gd8r9dY229vspCN4RpRb+
7iO+uj293SEhaqrEQPR2FAVe+cApG4/DVU/EbhGxzWko5MFE30BBE8WWYlIAQIbl
xFMLFhojn/KSbIiQK50WwbEojJOx9N62Ygswbyjz7dELTiuyBwHwfR+obbQ5deQH
a+AnZ3T1iEk6Ukxnxn130m8sMpBKBL0GPissbh9KqWvAkTXuOW7Z7FUtZRT2vCrT
dPwWKJtg/T/Ol8F70iw1ikbOv1QUUG81OOCfdIRKFB/aS0mlZTVm1iSMaFIup4+O
RqeNlyyOdHU0aJHr4wsVLdwVyRIorZEcz/kPAIsoPEn2khYgmglP/z9G5BNG5ImB
lUa5R+nyE+MkA2ml0KvqqYiFYA+orIBVd1aiubvnATJxQ8ym5HyFs9PGNg8h3lGD
u1CY8WPiJVzqSxckO9o0sO2NHajcXgRlnhHYzpm4C3AoM4aG/T4tL+GrPa9Xx8XQ
OwWuHxZdj3J0q0S6fCSpDjX78wbk1Nwpc34F3Ho1ln7G/fvTkp4WvkY15Z/HSTpA
D/0JokUf3Fe91uErw5oj35nNbwgzSynQVcZUHNwZMUvBxqw4T5Tqv0/1kKcGDPU4
F+Un7n+Za8wFgPy6T+wzKY8B0jFHWrruqSeBRBuIxzT1SwH0T+50AnXGRUNbGOZH
j9l489/8rFoH4pILvPssPLGvH4Hj9Ich2vrV8zlnPzeTi5e3ekA47QydpEVXrlz6
hPVyhyLYDcvnAPy9hk2iIG4nKg7/9X63pBPtPpih/ZJt98OQ2z9KTfmOrtrpfDYF
oaaj3vdDy55oMBwd9Wocg1AIUe8HHIeu2K5/E4yK0CaQ3CCZ343evH7p10FXGioE
DLGWIJqCQYaBrIXcch3RNfVLLIMdJ2H38X7Riczlh4i1AgykzhSueO/7Hm2VbFzo
+hT1LLq0XnZtmYGwUea5jTqRUzur67E5YgoWs0XDI7Sf21Nr7efAML7grCPtgeXH
uAhrEHAvELdCrm6OIIPd+NkGdOuW96u6eHFyqwbocvrpHSUaEph7DGIrHinP/ips
C0hHKZ1iosc4ie6vTzin+DMJ6FtvnyCGDkyr/4mIapLeClHL9ITpL06ckdnljuzn
BsfX5wjLhFI8NnPHLnozerCfH1wOnVYnYx8P9QZuNHzMiB2R8dAc39ItXTNFO9nA
QzUO1b6H07X5lqb+W0MOzQLSSdlgChyD7DJSfwFG1Of2IljCxd9cGhj6MTPGTybC
mPSRpEEu5M+hhBv6pOMcFMKTl2yI/tY2O32nlvSsXcs7SdFkqBZZ5LsgBLwXQoT9
LklarvJLGHWqOjukgGpJndTDrkEDsmjmVPTkdU1wiA4TwYIfhOa6euCmEc5dYRAV
MCnyBsUYTKeEohTJ2JA7Tr1I6cJCWBNIIzmlI7H/jmiMPC5jq2CT4JRyVrPEzS8M
EDSOYoqMKNeCy3b4skgVAciuGziQjUU1Qlbd2a0urdmDZSs9pGbZwwE0D2NbpICj
bIBORkS9YrNEC7ltutHrZQSZewCMvtE1d4KNp1uqt41LFJD2w2kUsEwPoNgYHbcR
1ZHoxvoZxxRRNoqaX6tb2WHquKFmntPvLvOlPpKEjMYleaB27gWlT7noCQFk88Fc
1s1+IuUwlB9ZjXwQlY11SpyMr8Jw6oPNPWoUiRTC3HnREGVUb1aXKath03/YypmM
i49atmZe1irtpxu8yOrwIvLaaq+dGF1yLr1tYo5xh0Sv+5oH6LI6aTu7jU+z9MnE
XLr1jeqIdLUXylm+4wGE/4CY8lYUGoEENutX+DReF0HYfLYF/TeuFW73dS3S3R8n
KrdES/X3jxDJ/j5ozqhpdLf/HLk1fXtuvlA/R+hXT9/l3+ntqPSo+hu56uYpPrYZ
0Eo4+AVAE9xvmjfIQJ7mCgaU1mdZo5WL9GIIC2Dq2eXPtJ4o2d9/tfckXd4YVMnx
UsPIs2ysZcRMLSTrMMF8v/vSCpWBcrqWq1sl6RCb38QFVAcDGqt3gTeVTY+SCunc
xN6fyTsD09wV++WFuvZMAYu7AUiBIxgWVOB5XTQ6heMGi8v6drhSSHxsEMazobBi
xHYV9EHon0mLl0jDgRgXT2YveLksl2VUMumLt4lyaDGbDYfXfFZBenfcpHH7anDD
IUFc9O7Q84ZmIpbRoU2qOnTnell5rMYEDDQ/V/Q3nqTNl5qhbZLuNP9RKU3Rxvhc
sry6XF76kasFDh5YNBLzFzs1nDhnQ1+C1YBiGfdpBlhHlGNmJ/DzGVur07V6OZxN
rF/mR5NXD8qykQnXlTTLTe8fd1UzuRpbHw8XxWcM/sBbiJ8la0/Gq5Jd8XIK7Ryj
FT0KXvbyeTfm5eQFVYbABLRlPJ+WgCGhvwFDrLn1lTwwLTr2p71D5+bZtmfjd6hI
qIIcYfi8uYiXhR5akaoAQQaLC4pNzGV6P7icNY9tQWt+ySj5Pbm2J4pgQxdPpR3q
CllUfRtaXU79FkdzgU/me2Bc6AO09jKUCA6NB7GVNK4Mna8zcpNQab3yMdWxIn+1
Jo3JAy3q3GfM3sfU2yLpa2BT6iEC69p0fuS3KxkRC7l6mMwAofhmpKjnGMT+dMMd
cZ1fmKRNlzCRldclrIO6uD3hEyNQASuLiSwD0LIg7OqfsejTbtVmnSKlj8/M2ZRI
uveNGMRNEodMm5KIG4x4ENJaiyHF/Qbvnzj9An5ipaZJnhIR1wn+CCnFs/9kf7T6
dgQZ90pRbBdWDTnBgwkEXM4aaFZUwgrm63Zntiy0toALGrQje5yozf2TvwyCsoL4
k0lYxB0xNakbv1XQCp2PM3iG8Q9xbFfNahG72of2L/2n7qO0R0NckDpc/Oyjs/XL
MhHeYL63RflBfBJWCs6SSSb7Rr/Tcp0sj2tCx+ilQj7RY0nTfD2t0EqF/EpJYjzO
hfcbOlYxGTOV2ggZTYNKabJIYYMnTH9yeKaMQrdO0tCWkN8dVv8C5I3hmVUQVVn+
UCt7KYF2ojY3lHDrGZot/kGJNnu+oL/95Zo5/bsuz7LTPMD1d2AMUeGHsuyKKxe9
b1aTjFu9/HTEAJdf+Z+owa9Ezj7acmAdklBoYHQoiySLuBDwaaeG72C0dvhDI7G4
D1QWv/ZAO+JJsUP/9BsAjKEfBniDalPc4db6U8dOnRos+kSEVXoaMKXVNEwFr68t
u9CWMb0eszoA3+UbRNwA4OOW3yGkF22TGCbMnjpRQtVkdBVvBp/zA7tuOusK9ZKl
czk/sBLQyiSp9pskyV0Wrlt9y+T4Ul+08WdY4HeZJ6lpOMrVJ5Tjm6LiGDAD0hoQ
ZZzn3U0YI6LHyoEey/ZC74LsuyrcKZd5b+lG45WwhDFi2JDuoQOg0DAcu6T+JASG
Hu9j1Q7ZK6bbQcBTRGOsYvQ1N+oGFhHhwfawhQic5PItCznx6GN3zN1i0ckmARsl
jC1sPYcu0drfRp4XXJLzll7A2OeaGel6IrfTa26P3Ii1Tg4GvsRquWPsiGGtxD97
os+fUWRAYlxY1f68socbzuN3xaOz0Ri/LcL0gpMYSinm+wqF+xoAKshnRbQLdfbU
A4poWcsAJj9Lrn6l7tgcVp8vXxtFsMkaiPvi/4XqW/VMI/9AFeb2d5vuCuxTTDdf
ezPvUV+bMnRp0BFlCsLbjjp3uQa/jZ4gxTIY9yf4PJ4SOWgwB+j8szc5m2rA3ZVn
J04PTkqOe1iCZIbbM5M/6v56QNgcMeKuYdM48GFIS6Qx5WhzylOpcxbGnmOhzacT
aiZL+wCIfNZfOyVX6NaayCi+df9ZqUn2XPRtKMoEVBPUIw3NZZdzgKbGNcA0jfak
PCVqQuR971emPlpapPIDlx8Otp0MGuNVdwBJbFDfgaLFWpmGvGQr7PmmdilCKxJo
2KLXD9rtvDrlv1CRNdsI26YQP0HONxc4/dg1D5vMZmu9lgZzp9tfc4HVwpN4P8t2
hLYH62/fIc4M4peWdGehpzjxL/5FN3fWYImTOvn9kQT+A+E3iuEM95oi5MAc+d54
ZhHTx9VSyoFlbDbVMwaFprk7JOlgUgR1EWtjpwtcSeODQQqrOoLmphkPmm6dd/BO
SKlKgkSwuYcm4pcud+lr7+aplKuQxrff9NsAg9GcdYe/DOR1e4xNXv6YAVsvh9en
UNVI06YCGNpKtytvFNtv3TwlvrUmXLzEYCyezOAte9o2Qy94ldVvDJG8W0yDHqeN
XVQ8TLCOHSkEVInfMytoUifuLpr7LS6CMuvd3t2SKfFpHLB9zOeUvYDTxCsiXNmn
1rufBqHdqfdmS0sOgIdSaEBQT94Cxiy7uK5kAWW3xz53KxBY8NA2X3wIbeRR13ay
IPGc/FCZIlB9tgP/RRLHZC5ZdqbX6rB5zhfgvPWHXbO2THA6/hAnAQT0q9rCZsou
WxRJLEndRR/+ATYI5ZRWZPr5TZWaMkJcJyyjXIeJPkzfojK1sI8k2n+8daF+Czok
LVTeG6f82Q23Q67WkBKGSumop52K4sdYnDSbbELR0tQPOHo90WLwrbE00x06tkdM
fGkdaKTRyPlXuZiVX4xhVrvMLDehOL9ZmrNBHr8nvaFVnS9CI4/ctH2mYXNWZcw1
/jQWG0xAAteH6AJ3H7N0pZFCDn56YG185hh+J3fvj2SHEHW0HBhwCIV4HqInJcmF
DjVJ0ADqe6cpfCkjcgig3sQgSgS11W8AL2s/OhGx/AVvPOvlp1JRoqETL6xwP3Q3
UnksEmNORlKEG+wOWUC8Jx7SCq7zS2QsMf1NyFjygOMzxcYP9p8H3zxaw9hBuniW
RaDEL2OUCMbL5pZwUUT3ack+cD3K5XpV/2kDIZwu417JUd5DAfrI9Ax5aCrdQ3FG
H/ODhOA5ShcNX9TayI1gZxS5LvQSfKNnWf5kxnvTowu6se4okqy2zPWfrwtp/FRG
kACICegQchrvLSc2AMtq/++HKIYgP3f63TeXPAuyzAEuz15K22jMGTyu7AH3Fcyx
e+MSzN8DUdwzlmadce2kzn6BWFQ/2kOO7C9noz6jMeeQE3tBR7gRN0Ytp1n/7Gkq
N64ITQRVR70DIJOx9GbzN14PlbpA8sLbOCN7fRDkan9D3IuiHXuWRO2G/sj7vgrY
XNjUKcylEeNSO9lKHz7ckaAuUzrDCTOSagpdDwBl0y4KsBiC3KgksWLz0QZcrCnz
3fSmGFzKNNr3TIBHQyCmMmGDUMlGrUUXGsE226li6oVErMaDkimZCnaXx9fRjP+G
/yW+0os7fPN5eTw9pkWJiolrlif969hlWVehR/VeXSDNdPCMmYAV3o0w5J+hSlLK
EB+aWrvOuTftwk5bQpj8fBURpVlahiJnv8S7i6LruNcdCj/KSZ7y1JJERx/Ryug4
sOXY6uApBl2vVyf1hEA8byUeScRfqNvekd1MxrMYWQ7aUuGRfr3h3XheIyQT2WQC
7kh6b/CJXZFcpquEjkdXKVJKb2mD+hCph2SA34SnhUcLw/UwTjwV44WR42uRuGOS
pSKezDjF4uvAWNIOfwWQvhrdPeJRnLmU3Bc5BbztjPtlodWfyRcVo0NblrlAF2Ye
k01cgAgo+4ucm/VL2Homsoq9/hfUF12EutaQHSiyhw0G/t65X6dapNkSczlRkOaL
vxbrGQjKTYsyF1bk/WCv6Gp/f015VimMnNL1c1qdhlIo8PWdc91dR3yKWm+v3ByN
bofBLsrh4qUmIFtxQZAdHFXc4Lm05NQ50caNFaJRQ36S1VSBQqGxgn+b7EO6Wgqx
n5Jnt9oSuHkF6DJpvWoCThv/V+bXr/3w0Lwh/4xLLtLPhnEWi19yJj5SPI7SEPKY
pKl7jvDNq6G++Yh8O58C6RwujYyziZKu14qJGQkXOWfrf+zVNWpO7Tb6yxWg7S/0
C2T9OB8Zvaf6QcVIgBHlP7Ad8gXH8Uo3M7CD6ywYpJMtY/UWtA/E49eCfKJ6nPQ/
cdJkp0MIZNmaNVa7UMljPJ2R2UoNmgR55Om+GcGcbh8dMCK4/iR2I/jW71iSrhx3
zzEvviIEId9S1AfIWX5wCqicDi1GkRmVOpS5b7REXEDnTM2kF8VGhWMoe3A7Xzqa
DVmLQjEzp0R57twBr6Q5KsgaVlTMCekRxA/wnyjtbLbbamhutTXKrmTxZj5Yw03N
D13DM9tuhkl1tEERjNHJbFGlPkLkyHkj93ZaBb+6Jm6ONw6RtV/J7MmtQbe5Ubw4
kgH065JJb3E6gwNuYoLaiT+IZptrEjvJPbxXvy+qB4LgM+oOWWTJF/SUv9mUbH6m
+ycK3z5fE50tPzmNnQ30MCHySj0tSAosbJT1mP7H/+Eflb6/Af+tkOF59JpSqm8B
SHXqhJWST5L6yTCLm8Yb4sxdjtOy2bl38UvRS+ApTB7weWAv2TZlrPRsG119v4CP
EVXidUWLmHrB1Rv3CGP715z/6BIGsZXa99NvhoYum59FT6KggzjVtJRGcMse1ilh
zZYKFmx2Ea1IRrvM4cmffiXorPq0EQ/3i+NCvUWSpjUr0HZ+BNg/DJD3YEv7+UuN
6+khxqYg7a/d6mr9QbENKUt9P1HYeO7tKbgVjMXW95q6TX/ER7WdyGu3rqsdt3B6
UTrxpsSlZcPYltsYbxyNHp2RSHLPmG+02yXr18mSrgRmsJKjr4f7VJKjmKMVMCq9
5eN0XrCtJPoCI+gaassNR6Yd+vtfzNEE31XfCjUHdYrCUTPdcO+xELN1FE+l/Mr8
CDZ6Vc+1CkEtNIPD0Gtx4uX869bn8IBGg0aNhYhkBAK402DyE/4XP/Ffa/RR11Eq
y7yY9nnIdHPoHkOkewbJxLp1YQuy/KJOQ87itAXuwaPbFSO+c/BwkqjbSswk90WJ
N025Z4gsV0rxoyEld0b7USdqGsJk8mSNV1N7ORZelZKG7r3W9bonwfP5gIwb9X1i
Pnl+V6udtIv6Fw4olf0RVM30EbP7OPaGBH0d2LegRb3b4qMI6lGrcUiABL6EtCEn
0CRfquCv/ktdsTWnrrV6Woqcos9balADfdv6dNnaU83zP/is21iUNWpSdxV3QjtO
TRTQ6IXRnGZzk0R2h6L27Gp3RbQxF33XqWCZrXOnMBVN12nPG8epfd7LKsjhzq6d
iHy3Xa92eiCAY5IpYws2u1R3oYgV/GjbqYNODn5FW+1wlXAWz2m2OdiLrSjeFBiX
hDe6NEjQpPaOH7xHOsRqWWev3LZ1znhAR8DZg3GxFA84o87NryjZvaK9AocLFlFO
AyqRVbbRKnHOD9ItyRWxPLmQYLqLn4A1wqmKFvaq7EFBOdPIjfw7IcjDzUHgI3s/
cMuXDjAzWxEq7ZD4aT3jaIMuHZn2wfXnpKjVO1EuN1AAjFiUtjWTMOHs2xswSKCd
858b16I0vhwZsm97BrEJFyxYKdBkX0NyQ4byNYv4m8fIyNfUrX/KFzFD1379XKZn
+BM2UGq4oU3emDgFTN9VNexLAmk2s3gXuIsUqbkyt5S+B5XU9qVGfBYZBkWft4Qt
vt86BjsBPzxEj7YTfroMEqRtNS5AggobpqsfJE/8HUPN+wC+aDdRAoUOTi9OANtf
zEbrxJysWA16M73L+oqlQ3hRmxvhHGyuNfVD4SyBYPKRwi8J83h5UObCIsov+xUk
prFl6w15kkCBlTYi78jKtpfrMipk+u2UDhscAC7CjZ0P9ufCgPP8Bykgtx/xjEuE
QPVs41WCc5xF2ak+d0e1x3b2716gmyxDQysqPj/fTTJI9Vpj+u5ixI1sYGUvdOEt
OnYoSI+/6sv+nStgD14hM0yZ5jFCqosZGuVKJYcnWLFeN6SxtWrU+6Seylyd92Az
hnkmzt55LsFUG6AWbeRLG8KF+9k/zKPCEW6UiU9XtbIYYlEvx2RIlUA+CUoTQjhk
7Vj0rL5RKNkUcGmNpNOa0izfpJY5mrzRB7UCH2/LA3kVFPP+D7+3XNnqIlfuYFcB
AfgCM5KHHsWu9wCfNPMdyqlcvD/TKsVPrxiJeAqWo1ff0xJ0f1WwSYdXE0d78vUi
h9K1sRtkCRMkFzAkXGA5ZBKyywx4i3ZYPhQCSH+g+q6wuMujAiaMJbRnHwF4Z3Xn
l3V9ZDNhf+0K4gT3antqsb+55dCIDqTIDDnBmBSbFVUVyd/uj5SgoDksxMlXnAWz
8Z4TzxfZYkzP587OrqH63/ChjF+1ivg3USeUP2T4qDruLXhvrQ7k0zncth2/c9zk
QMZIQx6s+baYMf0eavRcYTaZVoeyx3p8Lp98jO8g9Ux571g/0ah8dESINIa8rkSw
c0sEexbzfIw7P8zETe3rsOCRJIxxRZUSbr8LrYMMf08+P4uA5sRZ4IYS2RPM0JXO
qUBwAFjcT7VuF0PKrDT7Sk8VdjP4oE9/vO55ALSk9VSqoBlWZ6uZY6DSr1hZfvaW
9W626nNM6eKbeQnuZ9npJm4FovQIrJNCeKHnIcJR4zyxXzEad+Q0LHmJ5/0Syjd9
VONcZH4kP044wHi9GoDTZsam1vVUw5DOiGTIENR4XEgbRRi/GqT+hP2qc2cGqOGe
w3ZddRtS94lQVT4BVfc8el3xFd6f1mpn1qZ1rOimezmfdA2f+AGvQMza0QpZlz7e
8voNShFmeQnZ8wfo+DHYUnmsQaYf3ENwXX8RdwT0ERAOSMZLEfvSN1uf539Sug7K
z8gii66IvMO3JtYwgLyNTq535mGjp/3jAG8a2PJWbL3BffARBjSDW5XaBOWucHqA
JxOXqTFKf27r+yYKXaHnglol+ThwmXuEulPKGdvBwtT+qHHt/ja0qBywqgw7EDqJ
4jSaU/dpmWBRNruh7rOF0lDtyEleAT0D6q7KphRH+P2DlR22vY427XSS8nzZ8PUE
FgRUyCCz/7RQZny4exBFQKXpo1/7xPkx70aB6xFhP4FxEh5wcVNZ1EGG1/PsLjee
aSuaLW1GNStwj7fT5bptekoOhxs55vv+Pd8yCPewbUCKgdfPSOVgFpg+3IkGqs49
1qBevd9NWw+c3el3aPi0aKwffpyqGjp/NkJ9OE3IfohugWzTkXGabs/RzPT1L2Tv
L0KYBC7417XIffKs6jvuqWih2rTsZEQbiLRWrq35kP2Tf97Y8QYtbg0DqrybpaKk
fsBCcaNlPs0wo2Gnq1NMvlkMtsypH/9VKLdA8TJkFcid3gRYeaDAmq0U9lj7eB10
RDz+TlGF/4Qi1u+EEAL9PhMMXvjHPhaC9F3JFZ5ivCntz47TxairgUAqSO7mjjte
F+P2kzlQNEobMajwAml+UQyl6Wqs6yOrMLdeoCqh6w+UlUFSY3q7GiSLmDMm8RjI
Omep14uvO4tBZNHvU2S4VqwZUxzUgxVZKz+btvJxK7PykyVuuPHidhisOkDoyUbi
G7DmbIDnuVk8fwKl5DHmluN/F1njY6jF5Af4D2FojfdwjbrVaRfrlcbaPiIDedsL
toXBmpTTXqcebcDh8Wo+SXgG1H59jFjNYRertTC3RbC8gkEBymwd+V0TrYkz5zoS
Fjd0ep4GrADwczRAxKIbhjhQA48Ze6blikXBA1KWTiv5t20RJ1gdHgqjrW3h57+n
wT39I7YSbjHGlmstG0ACcelvNtUG7G8Sj71KC0eSFwP8jZpTAzhaNWBoEMtb4X0/
ftL562nz1HojtXxmcvpC4tgfCRc1Qz330Ie2Y0v5LZ3CikD1au1+7iwYHF9nYhm4
cLJl5tlY9RM9DUd/EaBakSq0OwhHXHgOdzb8xC9uA6a041e4WFNevr8VmHbpBGnQ
3mrhAqZKh5hg6vhI1XyI8DKPOg2d9B/m7OKGQgzIpuDWUvFqCodhyVwT3oXVXzee
yObOKXeXsxltmxkMgsZPvFqwhfeRTrx31BiQDbrdirRnDu079VLGNkk6XOgxZAPe
JnDQU4SwzJXibwx/OZBSXtkXcnQX2yrjs1t52+ZBh9EyNwnChp9RLQ8rXwgFZUj/
3++VGYq63SK0tv7s5i4UFg/UgpB1NpOdPFRNRuVb3gfFmggLTJeHu6zvg33du/2L
yPoFXDt1gc8DAGyahDVqtUdXf0jmTvp/8lNvs9Xbn7yf4BMyJXa18uYKsIrxTGvJ
iHpc+gklxg80dGC2smg141d0J5rmA0tgYMcSlAeZvZWgHdyieIMeNFnWoA0Lqeb7
Stay4SOQGdgRvHwijiJrMWJ6NCsvvYivWbUz+2b3vJMycjSQRjJ0+nZ9qcOqEiub
BXDg5KhvY212WnzLkLtzMDBsPA3e7fytzgw67fPjgwnWvhNJTFAyh4vpYzsooSwY
pplGJavoKN8K+o059UlOloEVhnRQ5pgs3CPmOFUOfAoOcOGGq8Ro5iYpldc08aDz
PBkleyfIc25LGjvjEhzWlVyrjRuFeC+BkyloqU6Fsiyqd90EG9/wGXq636w1a1AR
1AWZLM7o43HP2nbcAUUswZukRDM/7chVg5bqe0FxuXdmoPvX/jIISMlWtme+yYWC
EFwEHa5aCtmer0FOeHboxPgxnUe37i+ZPS7UvcFWLx2egGUNtctWDQgOssVvCO4U
H6Zq4hxGr2J9IXT9ZrKv7jTON0vSLdVzx3TYg8saxKYJXiETU22ZpCmhfFuDv0XV
10RR5VE4EPicu7IyKie2hG5LxrktBHksltgtg7VhCplw2LuQ6UpeKW3KbpYWip2g
yduys98NvaxrBUbHQrVQqMFxxmXV/hK0twXBVrlal46ldp2lJMeX0upSoyMHR2fm
UQjPVCdnJQJbHy8WFfWvZGulhucdVb8xN+dKlJD9VL8AQCwRAhnsyhjc0WNedz9H
u84EsvT+7vU/ICMuogA8pLpz4nzqyWk0Y56SSC0g7ZwgaR4kvcBYfZ3FeaybAMuU
sWQK767RkpeWC/5lsghZQXUsujSBs/okWeozEuar2ZcEbI5+4Y0zX+LisdGKM/Co
ENphvAL7irICMuRSSdjy3/bZK9rnXpQG28IgKvS8TenUxIaHZU0BUIlKMUB1lNyK
NHSNt+TD+5tyXjooto62RSH+qjGB2lh6XbrPptIW7tQE7kB6jnQ+TKTjMvU4do1V
18HrPMMOChVxOouVwgxmSkojylBXAYBJHqgWdAjrd2C8W6UbXem1WUDgeRDqPDs8
JRNunaLKAqWsLlSM/+uEJUEC4fbB7lKnU+vxFfS89ol7ArED06U6eH5Gzd7A/6WR
Gl+UKD8k2iaVrvQKpw3frAM0F8xyVpCWSREeCD+9HIG1uc0cG4KtWJcDsxICWTE8
xXBdI2b8tqJ6qhAOhdidBTCDPWJfcmATbT9AVY3e/BqBqhhRaboWxGIUCh/wvJop
gSR9hZUkH/vkvp454Mgod0lup7+biX9NP7ualpJ0Y3SoXqCjmc+jjFCMe/2Fqcg0
+P1Cfh0HR3WNa/s1NSMprsjtfcNDv+n6d4Nya68Bj/OgeGVnbrQsE8+GEnoANv7l
Hhw1Q5GEcfkXQ3z+Z2TPDQV/a+A3MuTFV4rh9/cAV3NUCo4QvqEvB0GljMVykRg5
oHfOWQnJKOxAvCsPwdhz5BiTNbtedeMlpHKSkfsb3648gG56P+OnSakcD49dLgYQ
cYNu9NgZkNeoiupF4n+BaJ2falDi+2Ml8AzBMjsCaZq/vIOrMkpWoCil3uBJMRNs
2tIhzbllqpP5rNwmI6lHQju9Y5L+jzE9KCUuaWH2yCSMYjgtoFj2OljwcQj0un8n
tAILEmCESirNMdxYF3vT8/yLxMPHNWK39aYYnk0Rpn2d0y+Eh0CNFbXAeTUhhjy6
dzQ8rLeq6cH9NjmUHO09SMPKwJmk286ifeuIqA3VeYyLMfOPXAloZ8fnQi/WcS8W
O3EwtBshL5qna6Q2hhMaWoK2ZFVZUrhHqnjlZGGrgWn0pH9vHrgP3a90ezf0665E
HGCTAxm38zNdgaRUnvHPVjy1FhWNwHA3Jo3+0C3BonApWCz6WFPySiihYULSXJcf
T0OYHQqS4kOnIDpuZU61H3fIXSvj+OabxEzd/aXg4RWZZ8C0zTtOftQE0ME0lb59
H14T0Ru5mvyKJ9RsTDupMhrJRcgR+atfFcxiNYhyKLRozQEIst2YKNL3qTmhKA5e
CrYRdAl2weRp3auRZTZldVdXYFzUHwy26pERqlsTnQOPa8sy6bpgujvELobFkdkX
enFbHwcrO+cJ1ea88scXOhvnp/0t540PwbgnFNSYBGaarjCrg3fdRdpPI5P++Tld
aFBj2KRuT1VYdxihWtQ3KKfXzGEajJSKjqOn7zAk2piRKtEzd+qdtQMD2XfvEvk8
zjRPo94TNqve3eEgE29V65QGmhbetM1kck5A3XtgKgIkrCil2ZWtsqXZH/LdOkTh
LzhO/D0UEjDdWyFUstzlB8bZw/JkeVIqnmirA1AUWINHIw+Eo7gP/yiqvWXXUKy7
4e+RsHV6fRhzLR9y+cD9x9uEu/VaAnlCA+5u6gpYIA6bmgFna6wYfUg7aHEzGCRG
1a/blgGQupMmFe9trHxQj2GeyEf5ORPq3aursQsOzoBO74Q6ZqJETJBSH9HdEKP3
Q1ZXKPCZgTmoqc/RIxZa4mUBz4wuq04cNGIg8G8V1Q9tI3HQ3c3h58ur/hhmkfnY
OuCwfPue+E4apyYAj5ODYdMQcaFhYXTLM4XSiaQ+hlNzTR3uwJWf4Vi9EurkHDCT
UzLkbGzJ8eo8Xnv4AYCZ3znis2Lo4+xTvb8VC7h/KvHzl8yCtoTN1dX6jIjZjLHC
LjnTop2aN4jKVjJPaSPFDEVR2d7+d4DyfiWV+HsGoeR2PiT2Pr065dy79WU41Doj
qLIZ/5keeZ76Y7nIf5kBNF6lyyQme3ZD91VxoteBQSCogxL6LQEjYuKLdzc032V+
OXcQnT7Wa9OVxe8ubK4B9Vml1a0cHb6hDXZqy9GVu/Dq37ZiNgNRqBSgEXzkTZa7
sVuyK4/cP3v3RlPZsXitFFrZk9wpfzV3yWQylqIZ9BMqkCD+5UpyV48vV6ByzfMJ
kdZJW+VYLxbcu+m1XCX6mOs269/ou+vJ1mg/RyOHtR1rwvhS5hDNVzv+YjuMqyp5
VsOC8TKG0KaVJUM0cy6Y6BEU8dTyrny5XaBD8TICYE5DBXwZ7E/wFfMygs4HemBv
BpcYYUIpwkN0dyLPBcqryWqHlyiKcQHMHQrOuvPz/sSHip3qnKIYOI+F7UyHS9U4
lEcQiT2QbaL3Ulircr/8bZsUui3Bc0S3jRDVo7NxI3ie74N1va3FP8WWGj3EJXhU
a+KUMvtXjlqGlhZvFlHRRaLpH5Y/qBkFXxhvXfP7ZgmkGV0IZn4CAv9kY7EyxYPd
4v/Ux7oS8otZRc7JUgPH94+rHTbmmLUtGI7Q5ylB/8m5WjeIzvSCTED0XW3yAM+H
X/rETPVJcYMEdeZoYRNOpb0Ra/gJFwGxDQejYOobyHLsbxQg/3ccBqCmjgzxHwNE
Pg7uxGhjN5RpSkbv9vJDFWdwttG70dzxUqSj0SNTK8ZDKaZamYnTJA6Z/CmrTy9P
HWpyaMpw+adxyLNiasA+Uc6f0LWgtNLt69P8qiPX96WQ7vvb1kOw5LyUcSDiLbdI
m3mbCz9J8tvrDSZxAsrma1HH8uaBECX0G2wq88vJvxSlf0+HVCajzx/IPEemwSBn
ChBal3bB7lNpWSWcAVZOKcWthX6VhN0yLTgq5x11AKFUu9dhZ0gwGI+B+XJMxJa3
TKNS89BW34+nFYol1frhdiw4gW+FGKlMA8nDV3O5tmH5h1xJ9qi+SKlxKGcc6Y9T
u1h+oAtzoKWNgnbc1mU06VA60s28q4mEPM3S1HreZnsZApxALb2wy6eDV5Io23SO
wAWXJMCPt/YNI1ciERnvxuaUOR4rke+1KNJZhOy5FyZgtJ9rM08SUJIsDaa4/d9f
FboUBC3oCIqy/Gs0ZBfbF9efRkiRKxtMPajesJGSHDCld0FghE6/iVY+WQhMzVfm
bHhFBdgiw+XmZ5vaCvhGRCLVFF9vBYhcchzf2OG6Bb7AqvRKQ1tUEcLyA4StUxnR
NcPcN3y1/pWXrcQczFaTVxOvJlYBC3HWGmrP3y57S27C7g/WMsUNP+Y2annM9uwJ
qGUhZAd+Kyll7vmrdZQfEq3RFQBqiAXuO61XlZqpJhg3Nsj38qbuYZtFORPDzkTX
moN3fDIP952TCbe3HEn2poeFsp09QDp5ZOpJW1sCdS9kVAKPMtw6nbIxguw6AgbY
OvtbTAo5j4y7FoYDK/ndifFrQUy3jEWA0BuXmVxcjWBACNU2LDy/YqGSBpU08W5h
Ahfb9EEgjeN38dTTdo/swVVaP1Disf9H68ySZZ6y9CHqSWR6MWfW8DkRLRCfCdAS
dg4LtWYXvfRNfYcLjNywpCxAmeSvpJM5bhZkrlnQ6qQIU/u8+u4CDL/TKHFR5uzZ
ZlMwSZbxSagPynY3JrZHSJyTtqgD9Dch4p2pxZ81nQrusTLohKJsbzRsHbFu3U4W
ts06V/L3YZpQweTMIbDxfuzf3w0Fme+GqADOEfL1oEbRjB5WV9VSyj2vYVebHmwm
6LNtEK4waZ/I7msJxY6gQaAl2+1pqJDIibh2oqfzPkhlTh/KMkDci7DH5h8MFJ9x
iLnAHqC2eBNpkUxEJLIJPPJCnL88MJ2w9pD84+9nMiz8REAADambm42VisBv7LXn
8sZ/MoXbU16qJUIH6umwIGBs2Mc6lj654Aq/4dIEnb4exKJSYwpg4WtMBqZj24FK
uDlZIyjlbDT7S566owNCx/SMcXfljFM1Etd9Y4d5o4S7eHuhClbgGWNmSuCgRqgG
tSNC2AZR5KURRIiCv4X5iEpBmtBv/HqVs39zEB8yWMSZZ6gAncQcyyODWamSdY0K
QmUPUlSU3GNUE8b6EnaIfHV4KbNsVXGIcvyGu75WF/OK0/h/3Nu0DTdxVi9I7wo3
uaU3+WVnLa67+2aaEwNQPwNXaZw+3RSAa+9CD6a7XGPLr0YX2Zui+2b/mYuiYhfz
9SpsKQ0AGLydNhWa0ltVu9XcpYeQGtPuIFhHvrkY/6W1Q57QhzMPX330w7BIEv0b
WbJzDo6NtN35d8nM0ykHaY/+ok23daY8RUGvvu2Fe4eaVhXm6EEkdK3oxlscJ0Ug
z/Krlhz+DFnWXX5aVruS/mI21OVPA8tvIFsUklXApLnYFFuwZxsq0lLA/fMieV0E
JxOzvPK12jQjTjElgsfsnq8+Fsb5OVflH5fuSweHyMm7lo5demPWfA+Vs4p3Udnz
jflNHgo/Uezu4f16ewJnWQU2hSSDvaGs13EMHwMomhtfNVXK2+ACQmbt08WuA4tp
cTlv0wwvHffxwbj49rj7heyJ55vGMAnu4zZRv6TuUNmUYpbRBa3tGZ0oCHzzgwHM
PIKmBo7oXJBPDo0jZGwNXmTRabMJBjr4shNjK00E3eM2aokPy7V/b7bkIARU/jM7
kYMp/gdzDcst7ASrd4yD9rR9LTra1R99uumj+ENM8oV7p5NhMSOrNrN1u1uI4Uji
b8uTA+VakHTXNXvIKBR30Co0fafj8AtiT+k9jGMt76KFoYwLlOE0CHv6q/mPBLnJ
wCx113rOwX1WAQMBBmjGEl3tyk53sRXwO2/Gc/AiM13WHESipdE97+U7hbnCXSeE
TxI32jHM6VHpVtJLKdXyNfhZ/wntW9DO8L8gyKERg6xUvYpOrh0dOzuunL9pKSCh
+15+WPI1NJvkkOViap4dn7LV3Lh0RR3J5G5Kp/I3XNuqJVAPKuLkzbmUX+s3Et/r
B3Z4l7OuABTrXt09uGKVtHpAQDcmGCl/M52i93ArjvYWmJUROdAz3+TSgDDPmW18
zVzZr9omfd93dbkfLwep85dM/+rlJN8KRrfz+naLCjrE9e9F176oenVBSif2QGVC
Dux5xihUzMDNiPbQilI1My0clq5KVdzFZsxRWLzexC0+MVjVzkGy4I/wjFmJgCGV
72zZ33uvH3xpUCD5X54leYBldriu3G+8UnFXh9cFPDgbZcYyvrT/38+3a9kZR8ta
7yD12gkYhi57xxquQ3x5TVAQ4gIdui6MzvoTKW9n5JIv7A4uT08/PVJpxdAi4Cxi
3RIy0SfIlRgaIgf+kpwzEdBuv46qyDmOmonTO549bxenugL04JU1qHDAjs0bkO7P
R9qsJUQ0aQPzWPmmDFOff3zYOCcpdiJkMdCxW3USzOxMy42Tk48Nss0x7JO0viNA
NIlY0t/CcyT+RRuSGwHCC9RPYrqT4LWdgv9esS01ZaeRAYVJT7j+tvzjXtkWnjz0
klmy7T/0/PgrhdwVWsiLGqa0YACF2dTALNt56umadnFd6dXQfaVB1oM387z4jZug
DjdIWnvr/rb6feUkJe34iaWBUgqwHa5sri5FIYDYB3M53gVNnzWrrt5kVryLnu9x
mwbae6clxb7Az3FP3NpftZ9JFu1qD4vxFRt2f7Qdwe7BNY73t/h+mcgUL7+A7yum
D2+2006jfJQSSoL4k2CCYKOP8U8wm3ZN9LfXz1g/ZPfwtEVyX80VvQABi51ScF4t
UodfKO8lWPS3EzuD2N/0FA54kdUN2rvBLnb62lJuoCp+tTHQ3XYl/eFL04NoHKuc
vE8W6iFZ+ZdnTPQpd3td8qPlsUSaudc3vkC8f4DC+SV2Dh7KNBSNcKZA8LxVfH66
b0KriPkutLKRYV1Ynk9p7mAbuDcc5hVCzFLxYXVufOkkG/uVbbX4cvhOET8tgXJn
sLQxKLE6fIHxGScDgVNgZ3N/VJrd8Gamm9lpvyIckyyhOmbXFZz3Uawc3IwK5G2p
40qIKZe9ZT+EZwGhxPs3hr37vk8vYt7+xjcUSXWJJrrg8RAl2H6i/5FvmOLLWbjk
VNidlUrZnNOpdSx9gR1qGrt9j/+vz5QCoUfkJrbuUcNW1Qo0TVZbIW3K1Of41Qb1
QVTmhYREjIkdfDlFpJkUOPQ+rr5b1MP0heG5AMvuNVxi8WZ0BiBVoamCbunNZc+i
zcV2bq0Ui6o7aydSx6Bl2EzCoqZZN6IvXsngPj4NOc2PC5NjPY/EXGCIoYm9F9Rb
vJEI35YB/Y7EKvLh4e4tHOZCSJTNcbOXgvTpL7L4Z6+PAvyQeCzBJe0u+kUcL+sz
kaczmKyrDoY+IgPncIRfes6tHey4EhlAdriyet9c4IiOD6VFtaXF7AlnpkjUfgTc
xhhbBOdtWG91P2iVQUhlP/i/Wgh3iNdogyLAB9TAGTbbkrG9QlWV/BHkVFBbTFba
uvrdAVdUg1ciklg3MOFNCMYuR+/sLXYHpc26LvIdZeZh8ys+c+jfhPUyafC6Htaf
2ErRWCRmjhuy0Y76gTYRui+T/mNPBeh7m9QyDltMLyYYleMilzhAbqKfcswg3fxi
5I1fppZjky5PPcbX72HRcTxmSb+wwBa41VfPuLlY4jxF27x6Vwzth7NMWjip8zYf
SJCcTuQGMlZnGDK/7TaeLMKJKQxhLIU86o1iLtzOit0HwLSlY5AhFBuS2aFtQ+Zs
FoNTYve5Wx2RwCRkdwBWUY235Qile05FMN6cxOjJhQCg62AXJQPLDvokT1YOeVDW
WisRR21QgOVgH1hnuQBkSr7KjXlZ9B2Fmx4fJPthW5up/A9r6lAUI1HRHFzR5fmF
5dSY8jeOZH3cg0YZLVXkOX7bSRQOblteT7j1ShzzFsDhNggBBQ/A+0A/gJSyTgY0
YUg32JW+T44S0gxGP+iSLBsjFqEZ/dxqVqFVucpKufM72RQQaZQccMksVfxaoMOs
n+zsld+hYHa6qZrOxVoUFnsC7WlGPtmwKr057Fbe3fiiJ+xo64kJzyHU+WRlR0NR
iYRPt4uK2c5stwLzRcnNS9iANV65jnytmA/Bp6LhRWwLArPU+6w7FxVXeERGtlHf
7kZdd97ONCiG1577RjMq1f2jBedO3y5+VYi5DKVBjvhadYljj9hGjHNRPSPWUFWe
WN5e92MWbu/8TivCSxrrZ1zwjivweyvBDjn8q7yVUeGAmIzc9OeF0T/S9uJFqP7F
LkW2Tbr9G8HK7muU7STAmnwgCaPhNDv/gbe2j50+SLHhI5uEF/ouMKfPm17zYZgm
zipgVbcuNkPDHuSpbnXn3j6M3nPIfk25Y8rEHP5CntyaV11SFm8uRIQN7MDufTPY
DY1hlRjXchu5sWEKTQP58pcgdt0I7LEVuvjbTplU5GzEFz2SyuICc8UEczY06Iuz
YGTPBYjZi/T8YZVaJ7inwOytYIBFLaFr+pt4EOT5JZvW2CRVPB4cGfdw2xJth3oc
Zm22d8whapLZSbZfioUIEo58bVXqc34XxDFbv+zd7Qha6dqSYlYg+Cuq8+AV254L
1OrZBuKTOGLRpg0HjPzmhyIVsmooIka3dtn20dYE09OPkKuHvNUA2tWm7X1djRoh
Qca4n3CwGc4XGt0eiycL9Ch2+VMwL9pLxq9ZwVaoCB+IFq1ET22U8AjvwfckBYqo
k7MhR40fO2aYdajaQ5Osjb9HENH6Jygcsry3actF+Sr5HUclK61kVBXdI77eFD31
tunWUyT902RdbEDWYrtEXw2aN1//J79L+YTEHLAJyRIcZXBNBvzZsTpoH0T46AKd
LbZnb9sadiDjeikFkbp2Z2e64zvQu9VhMLcEsiMpvVdoKjCZ3LrBZuroGQh7Ucys
CMbhtRXMxyxkUvjJTFhO67zhu8cIPTGgBil2/bYAxsX92Pdp4IbDXcJ0OsmZORNm
n71PGuO2Y0/i567+0dq7r6KitbCqs3uFiUiunW1AX9M/B7VUw79bgU5rAznrI7O8
lh79TFeWW7y2M0/0fQEn0Xj2oPiDGEg9grzGlseJSn0rRnvoWRborBGIzSE68kvo
K4OtRJo/eg3ZZQMG6S7TH4CtVPXLwo9cVNRzgRdfMhTdxh44Ys5AQd/Szdih+8n1
G5B/Ettvfj2dl1rllDsQyHf43EgZH9qkpLciw4QN3gDowC7L954eYxo4a/DzSzSN
IlIwXAV1T1Arwy2hGYg9EIe11OEXIlmEHo6T4fJP7nhlFHTHAKu7K9Wz6hymWo91
jWTsyiH/XJ+dyDXN1Bhte4mIWoMWQbvP9ViUKHEu2UIaRQ0d55L0xRU7U7mDnbt+
ayjnGHPBTb4tkrx1KiG6dddGF6S//7z4iAmkRn9uyUkWGTvsDhwU/r3LVG5K1XnY
aicyhDMXr3guLUohDZxX0vbyBSRhmoYScjChN2iriM0wOqDyLr4XobYiDkqKkT7h
grhhhqpxk/GXZDQuhqjOEshPtgHu56mbEaaggIeYZT+0ocXWcVF5ka7lDI8vwGDt
JB/GNHyBhm1YtjGWKLMOm7vgGUUePGv55dSzkZXggMTiSiMTyz7DEEVGnK+Qnbbf
4obsar+jS/SRPczFh1UfV4W7dBUgZaHOTNJP+5I0zZFo+bed143tBkbXAuwJwiAZ
wUz/VKeaClmMOdgSyLbJofN4/FmcTWuY/pOVWKLnNtUAEKA1u6TaYfW84jrbaq3N
eE0j1+1mQx/5crLb5oqYCnSb3GL//ifVyNz1fcuk1nYmPF0EYH5wjGA68YwRaQPr
UnHC0jdyyebNosaOLwcl2cZrv4w+yZJkj6/VXvcvdkfIj/3Rcrc/aOm6h7WlNs5Z
xbrNiwjN8RMBmMn2uLrb45Y5CZhg2Z1o4U4v1m8ojX362Lq1h8NzJWC2s9ifIysc
xUP0RroaanJvY5P7cxHxV0D0LLGvMr4yYXLs2w1w7PiyPMvYLCI/9QuqLb77YmGE
Xdn8zEZ/7r/+E0+4/nux+Wj37xl6Fk5AYp908vpD9SF1IASKiCjRc/gK3N5YdFdb
JXyyNnk7dogiKlTjTqA51NomT2u48YlbLTcGaeTPWIydOJY4+j7SHABS8Nw5DJPz
FtOQ845X8XjlopE9ZUQy+tqz9IIIZgdS1kUYADBtLqtPd6VHN1SI7eZ0nL4bFE9O
tGO5zpbhYG9JbZkfhm//xlktwvo/u/rKlYlgEhikx4uYA39X/5/JFqxYdp7StTkx
wkJsVnHiJ9YYiX7dCFX/XJZujdBPLaHZ92+arcdmuPZ2axygBqC/43D1jEloZdpi
faI2TH7kYNiaAIt6MVSboJCmi/J7uYK/aqbX0mnzQCd3+rk1qUxr+ogL46Lsapsc
G0KzGO6wdrj7sbmPbrYzrJH2ZBmJU33HhdkNOsK7xGZHnSmZVxPjXSVqPdzO3BEX
9WKyKW0aoFvxVXTfv7I5GYkiOn0JXfvSzuQc2N1q3ya6YQ6oVJcU4hMPI50BPzEM
FSuhFPshGEj1lc76iN/S/MmjdZlnOkwDfDzitIe9gV9RMhsSXbUc8JYrQrV3g2Sr
quxrN1yzjCsg7kdtSfdw6mO37ETsUIMELM9QKX6F/XeBo8Apc5bnWcWwYVCzPV34
6BNfhmuzOISvw/UoqjDGW285s0Pf0ANCLZHXeo5fXUx/P4dYqG8Lhe2zbgQjI/NO
Y2NuKbLaikUd0HRm1LDnm6qJ705HIHh6weOpyp3pg6WP+WDvYp67xeSZHLRbFvcE
MQiQ2ie1tAL6T7gHoECzKc5rtffyjTmxQTdlDqOWtEOhxHhYRZXJSS9C7lxGkajI
G/E3pyN/eQv4GQdP9foS6QLNwsocVApHJkunoQERJtHj3L4oXWyZSNS+MUGJJqai
CGNT/D6Eh/9RZ8SGwMKFotau8nRbQnOyO9qTP80WYZhWbeXxVvoFzMCCUu/v78sw
Oykm6Xf1xLlpQa1PvAwnE2issmHgbFwhA6DY1TMUCKaOeHjgHYD73ppd8FwAy8wI
rDYQiZ1b+ShR1Sw3oav7wrL47OQ7Dx8RqMzEVYouV4U+hNAzm10+Jd/Q0lJkQ8CN
t0LtpCJATHdClEWpqqfFjr1G7IE8zPdykT538jTxSPryfy9gA6w6Hx7ArTuJZZcy
hISo5b0ZPSDGIc1RdMdY5hCjbGwgIJ3GMz+UUMm0AHSHMq11meSLCm0YWAjRHTLm
Pzx//V4oIZNw8yNGNEfjM/Up/jQOcAT4HuiE41VkuiJGqnudQ7t14yMoTYrGZDAi
WAcPhZDRux0ZovfOrKXdjd14hw2DAPrGsJBRX0gFqgnPw49irouaQlRxzIhLOLf2
8xvw4dQsZ5HiIvNT2NiMGAaNSMlV/sy5ZEBEjagLkE5+NOxdeBFpgtgUjb6qgT0V
H7yrdB4fhw3EQYLmgRfAXFa04ekMDGHBDznR++7FBwRz0S0Xah+OFQ1wVmSnUjZE
izpUvfOe8vSqcJhYgWpB21L6l15QM3n7iq1U/fMdUk8TmFSHi1cesY0avI9RUTQ9
ibiKPP/pzrR3p4HLm97Zc9gT6wi40jzqLlBEgCwjwnfy3G12g6aYYK7H16REftBw
Zhv8ctTpwsk5qnBxNIR2RKXEGM9kT3OtPrB/QGTe18kNvwbaogqxMDyKd05IWKyb
tMWOthiZG/HuJ/Db4ss8lOLpDDYn+Mvq2MxvOuExaRd2SQVT6OyxRN7SNnANdzX8
8DoJiy4Ch4tbRKQaM67F9VRUqYXWApYkj1s+3+ZnX54gUAVrKDmYb6Zudf7tjgwG
JsK+a9pfyo0kvGM4nLxWDcOxj+oHA9D9fe3Q0hbB59zxDRXGzdQoQxELHVVCvA6m
N4mJzl/3nW0nyguAw4EVa9Xak27xEYCWgjSuERp06yv+3CfFJ9lQyTNwceoMMNUq
7a7DFyJTuSrUs80th2w8lc6f+2kPKGcW3nhYLJI/ipmh6GyF2Jv6NR4VynJXhVva
iPTgUD2wSah0M1/pZZyn335xn9zZrquDMd0ksnfrC2gO8mn3I0bol3r4Twn1CWTs
xFTimw/RYJQY9gmC+bHfr5Ie3jxYE50awLx7WcOGxWYf86BXiIt7yoN3R0An7APs
S+a3pgPk4e9Qp3fwWVHZ3dc5EXlk5BM/ULFIdgTh5Fg9osQes7vV2+IpR0RpjynR
acLQ5OzUQxm/nILFUXBDXH0OtLB2wpEozwcrsH08mqWZl0RBFuCRtW5rWIhdF7vT
UTQ6Z3ETi54VbaNQIwoEezdUt68hV6rqS+S7b0avNWTLz0bh9XVK/2INfjB65d6K
6W0RK8gXJX08rr+5nW7OpaKYQaCtEhQaYq69O1NGzcVLvQKBKjm0tQHQZZjkTaDv
hNO089U9miofL2jMQqwpxS8S8rT3Cg5EamxD+jqzJ0C0s3/VxMVXwa3yQKYcj6Dq
zRPuB2MYUZX/NeeHB+wLs6kBafLwQ1oeZi/w1skPOiq2pLOY6JoihhlHGv5SMHzM
ldxo3xsdW1LgAWxyJDFrZNKcHoJnid3gPw4H7mWLvA86++senOar67UBlAokCo43
xDPT0wGgvFTSxDC9DZht/BebwJsoAOH5YjGl5OpvfZAibxXWzi0EMSL1VEx0UiKI
Jn/OKAl+n2frfv18YhBfexxWvXN0kT3gGOnDJweZQ5afQR3uERnKFRD7xXO1LpVa
+cKwue3rdkuDWvi+GYhs5tgXfj6InxTTi0z0OMr/777XoCKn41j6JMfqkBmLXisx
9Rp4o6vRaKNQePflzq+Bz1bLM1jYGvsAyt6m438roD6sN2xLRtkDI5ZJgvIrjqf3
HYaaac2WRLhL9j3wuYbAVb5IGF2Nq1FV8VnWfiyx6yYNCGRe7QedO6A36E5motkN
iB6yAH77rDrNZ+flgnei+Dvoyz4LRm71zIZVEi6pnhJIUtTqMspw39nrdVIBy3Hx
hWX2RcNyEI9nhgiVPjpboFaMUEvI5IV37xt4fp8uh7CbCgbRdo/5xJgsZvlN1tws
kTMyzCvNDHFXvIjJyM9tqvkgb4+3+8lyiD8YdUYYtYbQKTgu3XF7rg7he2cvg7y0
k9/lDWwhSq+hDUOai408PxxatkYCic4DrQmP62FiV2xSjSw9NZWoUaBPaqkt0Do5
dnaOq+/RETFh5KZH2Kozxd1jAo6THEf2UAF210Z7gJQVH0bQvJgF/6INwFWQ9DK5
DpN7Q3XF6HBt/3zZlnz23XrLirKOVVBVcSzRWcquzWjpEGH8hLm7n/+hAqWdWVlc
mAJyQ9/RxfCEBH9XqWuiWIMGzNF3UdYG71OVNycICAzvmhvKciUXgJsVZlDRAJTL
yLUJOMLw3RsWKlogsLW/0IsyEIzMHFrCY3b8mw0Gilr3luHV/Mseelh+vomzmgry
jL6uUV2WQ1d6NWHrU9+6ErLGWFcMg4vmOiYRpgG4pRV0NkxjQgZtseLvYQQHA3+I
Erk1femgb36AvQItCruhFq0m53TkloJmYcANCe6o16Pb3wgsMGBgeqIJVdqksDN2
AZ8nEHPmCXqhVtCTBK5usMCLvSFruEdY8ZRWaId3hWOmei0FpTb4pf82Vy2JkZg1
eQTZzE2Hg+wDFRCGNL+8sbHghyEN2aRNcZfmOeqNxxdz2cDLN4O8+glf6UkhQf0z
AdE5Q5FJK8UJENKjCLi1CRpHCf0FVu9TcTDJq0/5rNvU591U/nBJvqGwIPsGTZby
7+ecyeulZyzVHMimasUUHrfbHqn4fObRmlbAdK8OK+DcCMQ0Z66aJ5q1fS3UpMYf
b3qiC1HSknNiV6EfsIYiwZsmIgdWfObHAX//N2NF8cyWLW2AMYlQM2ZYW0JkrGye
AenEP+iiTASH0b9pZK/lhsG9BP6xrYq8llEw2a3/zmo++U8zs8sCBRNSkbQolKjD
sptYsOYOwRYEeYVNpHSlQ+XEoUrMGIdzq3dZyilzM+BNhcBQ4VHZTVHhpQ3Bjfox
wG7WwpQoZbytFuFsDsevQfgYXOOn917rFRBwpXorbAUrPTRwuyV07bwS4H/8Wv5G
5sXQTnTslKJ7t5mormsmAAQCekeRcKOzw7jgo99trwNs3DyGbZCWXXpv7nQHgtzL
G0Q/McNsl33moqq5gh2UX94UrCppkPi6dk9Y6yZEAW7q7vIdsBI8g8Yk2+dcsjJD
ZOsE0A1l9EgaU+S2bjXPeBVGUOEwJ50GgrTHCUSdzA1fOS8BuRW9UDJ/zOiUMbBD
w9hwBBuwCaXBsYw/CGqp+hXYS1Chzqy4eAHGJMubLZR6cALGTJuiCyERZ+WE93VC
3OjAOaB9SPa9SNpvhNr3iv4cDVb7twolbaTOz2D2hg6X8MWLH+8kXKMBx11AR64E
Mk4ix6oH/YfyljBVDknL9EU7blhnH1jiiXmtcHC0m3OtsarDfe8K6WiR9sFERBRo
uvaf2iLi9Tyj4vSb5UdFxIX8yiqfx7Pc+sLhJWaR6YuA2UkB48JQq+UyynGL35uY
k+sGYL0Ycr5o+JdmBCfQL2qgCW4O8Tf50kMZSgPWrjH22P+mrpa/qf/tx17b1vG7
+ZVcqbxRv1JB77CWn/bx098MLBectg1Yt5h7cs/JCT93uL266n/T27zAjyERw47d
I9zSTYYltuLADGXXn7PBoLDEE33Hp+e1BH8S58rt67DvkVuKJfDJB23Kf9EvmU28
8N1QvdwEQPhdlOA6I6zVIukqH7u6PTY+4MFeik4epQl+0drxHbiWny+OEg2egh0u
bZH9gh+0jHG9wgIFIVQPVTAylsOmbT41E2sCat/XycJEFhKFUF0YNVHYxo8Vin/A
PaWPlxbTa9sWLdkx1hJ69zuMFFo6qftlbOPfC8OulrH/LBErG6FOJisaxiiEWK7W
lWR3q/pD6UFEiivUDYec7rQUw9qjpDHcprMdjlvKCbdOIreYNC/YiboWNyjoZUCE
mjguj9m+pMf9uRBBefud7UX9LtPxqupTR5M8sg+vQSuCnc4isjNneo5EBGfmoWee
9cB8WjwiJtFRKAayihFt2GusbM6hMZ2JqHkZnedV3tMpS1ZTiB7pB41KvEudQfY/
GjHlSWWqEgwxgweNCzWPbAsdl4NldvlXINpxJ9IIEJ+NrWpMFj9qURSNp0s/mUTl
W6RT728pdI9WzzKVm/ekfA/MpSyGMDTa6g4jg3ISJYDljW06jhPU46uOfCZTISNk
R588rA8CjCb7Z3daQEh4VGnq348YWMeIsTMmlSI12O5dxS3se+gf0RRpchJEkAGf
EDHgQRG7VgYD1u9WpT50g1r4hk1NMjCFW4cQ2HVqieINhHdvEYxArlA0mHtuoJbv
rdKogPP3D6TWPzMROqt1T2KdOGMYZS6qdbTi38cUIm3CDS4+oxgFyP+p63JFfFvh
qDYX2ExpBF0TwQ3crGxxduGeoI0ofS70plSs9AGGlBjfLtPPUnBk/6O0b+R9kKP7
RLnlJUR2O7ROUZQj//JpMTOmeUoxfDeO6sGxlgIoAb5cMA0IouZnIOmIjVXoknvv
XOQYTo7tTlrlbWcecWYtjX7bui2uh1DOyv3Q9MoAWKkIXEAP1B+ML+Hr2lJywKN5
dmATIzSTdOjste4yrOpj6bijAc+sLy/rMwEENzjLT/RlAlnc1M5mrHaClWBkqegy
2GvePlLOq1ewV7l6AeoQ/sDJNys2mI+qDwBwcDfx5BqhUSfiohx2G8aAwW7PQKAn
jzKWhdKr9/6pIkSdzUG52LwU5smYHOc8POaZAVEYV73wFHCYIl5MrcvNUoqreIFL
KQd6whzzf0MnA9OJfZ+3Pb1om5d/7sc0auxbUUAQgfuYQf2ZIaiRJBG1atfaJEcP
FhDZAkDLbgFwGbKu8Dt2jTzO9SIQYY/WJDl7ZfBCI9ppWY3W7lcxpfyvPPujQbYm
0W7nJg2I393u3lsiyZS2aW8bxbQKMfI2pecX9pT4+/2AOp74/6D0zuXYjvL5tkon
SMmC24QJXEXPrkYQRdxI16eZhPoPOTAnYiUyl0JlS4U4nIiTeaMUC9DhhAtzTCqE
kTSnWN0MKmUA4AYrI3KCD77uZjotKAHkZU99FU3Be5MCTVcbOyqmJV0dNsmzcDQA
3Iv9x8eadg3/1mIlx0PUhRE43ZzQY7jUOakanbV3BoT3teqMZw7qV3JsWYGmyz37
qE9sV7A4LYelSCgjG6ApnmaGLuQt6xh74v0/RbQxcunnFWerByn1sECRipN/ZtdX
uPOdEjt2NJXMxSbdyXQndjo/M2EnX2RN/ngYQEANhPpikDoPc2WKqxQnYf9kcymm
yg02P385LG01/DltG6/EZNQ3VcFacFCA0DFU41tkhW7dWrC33oGORyR3G6TqgTYC
ChkwmB5Aosy6fKFxq+mrPS6hYz3TZvYqhEtQJcf5YykWuw3wtl/easSrRsDVe8OZ
irWX48luK6CE7L1qZO9O7TflkG4CnzY2t/tuKxVZkahubb3o9AOB8YBWPyEpiv99
ySNr6//QUM6LlEI16XAP8H258gCBexxDBSTupWb+jVfcN9rt8MpjxW4u4j1t//oD
lzWffU2jkCne2TWXOxZFzEXl/AghLJ3WfI6TrdL/8sgZRJ1iAULfFCoB1cId3jRH
7hfPIAgCAqxOOHac/h0T5qhRw5Rgi+MfdFHx0JIx65s6aliAGa994Y1ySOQxONuW
5nL5dbtm1WQEPBJ031XikmzscndSYImYiDL3Zh/7U5PLsrDHWtrPVJjzmejaH+ML
lfKrnsIOfv7x1+DYY3inBx8KGPdEg2Gn+SDKBeJFn368EE76Hh7SPAyRPjFY99ez
tDQiU3kbxKjeYiXsmQ1Zc4zDuS/q3t8jVU4zuhM81vprzl/gaZ3b79UgluzUBNpR
mZzZUGBkl26qap/o4KArZwgMcaI2IhR2oKWQHogrE7wA9qxu7dHpLvEbY+3GFdNf
Wf8f0X9d5jIWs9zqvIzcLG9OIO94oqm4p1CKkRnrJ8REVWjWttqkaKlLug6SRBhT
1+kbEU/xdkU6FAuxf9D+RgVQ/r/xrZEvN9AOb9vSLuH2kdVOYF6whyqTDcRSGbL1
flTrPYGvtaRLGl5ivfMwjWS7WsKGY77LiP0eSV+u1Bj6d5caWl5Dt6xR+VtsWd1p
n6v8E4leZlaHp7+aUnpRtOjCC9aGLWsKrnsxYagvGxHMNd/DjxeBfp73tpIbuqlG
ds8yHEQ6kP2QKwrcZuXF+5/FtZQ33tO3FEg7ecNkD/sezAvf06yUgRwI0kaRLvcS
m+PCa6xYXHQRTRAXzHIVxbxeOR0pyALK1eS+ASR7fHQ0RMEs3T298WRlzxdAM+eC
3fWSWqZxjP8L5HPVBuYnDRl5QjXeU3MWGPHZIKAFiR1OFoR4vg3g8BQFBlpJv+EK
J1bmBKhekJvFvPPhv3UAVgeEotwJzsS9FIBl0a0fA75gcMQUrPfkJuRyi5WDoyS8
9oz8p0y6pDrY6w9Q+1JBsA36+ImzjlSfo2tZbS6xZ4UqQTvxRA0fhI1jl4ernXlH
yzcvWY8x1lwDeHCfVR/ZbbnmuLu0bSsISVJsqlog6iovlv+2Hc1HtmwXQg6Eugdu
eU3XJROqRrcjTLA92PuFcI+7PHgr/WJDyD5cTq1bzhTAakRC1xNMuOm75qf5ea93
/cZGIDrcjkJHhlCfUL8KpEMS4dx/uEhj75TNdhobI6C5Ds+QmGNkut5RMTkqXJtU
apVtxem7n0g2A4bZXXbvjYfEkfhc8/w9MzJUqCW6iBst2SsrquAgBdx0azJbti1M
gK8IBOFVcfRbIJ5/NQCmAP4NsXXSaUoKimHe7bB8aU43JToW/UPBoZgwYAGQtrYE
IeU50T34UXJBL3UGe9RGSOp9c7QEFeWKzi7vGBTxL5vZcpT9MHc5TlzC2BRuiNk5
Ekq0Jb8n/ItqgF9K+6/HTLweIvBG6HcFU78eFSKH1Pdt5cOq70stUGQAIHZDkBHQ
IRABBOg1+V5iGJFUJptmn13JXolkrLi9uHLr8s9zMnRfTKJt8lBAFlhA0PWfA31H
Wn7cxTXAMqbXLlJZlE2GITySbXsUgzOCGWz0HaIlP83Kber6zRBq4zgsjAVMljyp
NDLoElobdW7t/+jhhfI2rxZA+rNZSbvVVK1ZAxyJyNSVs8E6EEfELltU6titbZEN
7D/pVwgrW/Y+naqCdHHkXILXcpkxY/ciXr058MSXgk1BBc17Y8iZdufgYTlEXqN5
doXwrg4lXWsH/xeX1TJk9DocLfkiCbg1TNuOB09imngTE+dUpJX0PnOCkc+ePFWM
QIVVA/acxHVOgPJN4pW66Oy57CloiIu8L5bbgVnlO2efp+0a6Y4CbKtvSU1gjPc1
8bCu2PEMViGxvR89yKpNjWRjqcX+/uG07PYKbhsgUIA/pXZ2+MDK6CuzT/kG8PaF
3f8v1LaCpSwXJX5DWNrQCB4UAqkirxDT61/7w13PkrmC3wD39N2FSdtLDtqXK8+i
uM8xVsGOtOveCx5PN3ZWvqIMxjOK9+JCLWDfIM8uahYBDZgvQzrMupHwQGhomsSg
C5MRtWssEX0is7J0jUzQDHXLcMaQXcP9DpXzHS772uglpAwBwZ/o4dhwUTzoh9hc
uLA5gV9LshwEvPeDidtF7U5per+rEXyq3dgzcyQh6zgg9CSxqfDYzNrlXOdBsq1C
41h3gCMXZR1MfYGvu1wPrVLFe33iGc9xg45WEIzWYDfJhJsDBY4KZ9HYZVpqreOp
EMl7QrqYHEjO1Q3b2vDxytVPJz0O5nN4HJUsC71XUDOyPmzBNOu/4CH2nPqmP3mp
Mv4uT0qzzXvYkSKauCx5LbJklYo0+YldGCjohHyphcX3xqC7hrpCgndbGpjrsebZ
e4x3ny3bqcC79qTDjpCeeP3NqvAsMMwU3IUtnVYbseIj++RGMoeiOwW0IDGxsCfF
ADT41LTSv2VTXvRej4Ov/aUKxEIijymg1U0tbj8AhLuejV9doYsd5laDTrzmniEg
K3HDTr4XnbX2aspJuHBFlqvKlY5rbD90cdxecUygnHDH2MG1Lx30pSzv7fs3Rd3P
Es8QFWa6ni7C7giRrgUx8MeAjAzf3Zmyy3Uq2eza2NOhkKYP0wzBtnlXaTN13wmy
lynOBubqVd1Ax38jeq1Ycg8qu/VezAALrqXc1XY8SDIk6Or7jkdH+HDp1iqS7SZg
ql3DLqFrgMHMy8nsVpei44YSED3/EuaA9NjbE6TXorYz6wUuy433mHORUZWpqz32
4lFnJ9fHX6j72sPrWZprLpnoHG/Cziy48y4pLcsqbFfmD03GFfbcJruSHydiCkD7
U2vVVvPJin9jWB0M0/MmUhSjAod4gu1U8dsfy2GN8dTTdRQzRq2CujUVzyI+a2+N
HhSLLi/g2Z3H1MlBKubFBTsL4Von37OoHEdcCWyD6yveEgoycj/KRU7moXkaCGX5
x8OLsifdop28j1rh0LQ6BUsCXqd30lzNjHDWYlzbSxD3KLNP+BJoxHS6kEykBOmp
WW8iGW481zTYX+6UnMcTHEp2ddPGD65Gd+N3swycO5XcXc1jeaxvJp7DBRFe/zwn
LbLYZmZqUSA5f62u3VWXROjjefe8I53JYdxtI5zO1VTvLMwHwZNBN0pFoRSFoJ9z
wepUpZMcJ2NPgm0C+zPeg/c3aztS2zc81LethVxoP5yGH5hbkK5qLUwYWc4iAqjO
Jc4ZbTNLG0FsJrPf7PNH1HYceDLdtru2Y6uacQjsT0urc/Xu4ttLnHSlZUXuEzCt
4ABBVLojNI07ID6485flmWSbwMpcf9VcImuuK2T3y+wdAtXDUP9hMcT/HsKfJetL
nmbm/ObIHbYzMsp0iuaiSHlhcFafovCvFFsmI2tonAXAZX67IOY6n/gmBMuinwph
MBpuu/23S8AxKKcmbQ1dpV5gs7WA96R7NoZVSBtrmb2rf4g97ccPE/7EXrdv+wpE
/B+/AdthArFI5yWwWVh3howSsTKbfPZmq9GDqjbJIDKpVXEevzl2+riOTPHQ4w+D
5S0rZ9GzGRZAcFAD9WY2TEYDeYgn6bnUEkgI/1mEIIKI0JJcmVMWZ8SAuPKA9rEx
H0HFBrrg3QS6lftl90+wUwRDg0Q4zt643HNwvdoI8zkVOpeQhldg2wWyGEjWP+j6
ozUQ6MJeBLswr0TvpsWQRqh7GJCpAiLqQRkjrSa8YumnG8QDme1uf2qHiApmdM6J
wzGgGuMNRjTy/gOf/MGUis7GjcDv2TIFLMuXoPjsgvAiZV0XHTmWTopwPWPrqXiV
gTcO6iQckD1mf/s44+Ab0ghBhPjNEhuZMNDU+yWaiEhN9+fyQPeV2iMWPb6v/48N
VsCsIv7M8uc3PnxwHmrWSD9aomzTfZB3MEqzi9Las30/E7pPk/zQ3oqbqMeTHenw
deo3k53gij2GjPgu5WIqJoylmptZEHrTh6JW4G23b28+Xetc1JNq5o9FI4at6trc
dfv+1S5hq8MM1C62G4kwIiIvr0n9w3UqxG/U/BSXmDa8yxTdFdW7QDkISQbVze0i
4fQny2VjXrsTdNDZtb7+/Zu/sRNmm7BeJvW2pRUGClvNLoHuBr0LMBpfhCPXIObb
mzJf0oxhvuOy4IToCqG08vkgSPO8NlhjM6xFbF0fz6FONyBaWP6GtrruzJbSuofo
bf04nq8ZTN+G2tnDhEi12twjRMWGCpiwc5NJwaEdN0eS6xci7OrRotgYlKd257E3
3XGTwWexuxKEgvyAloTm4IYYPr1bgMqghjAvIR3aYaigDSlKJvsWZ8e60pYsA5tJ
CTnX/Xkjt1lgBXvJJeXDgx+ar/jVm/W8ZQs+ID29YsQA6360OgxxvwR/yBPK96kh
fvMrKzsOxb5tG5qJeqjlhlGqB4AHiyM1l1MFjbkxJmLcF+D9zZs7xMUAHyoMWZ7T
F/7Vaum9MK7EL0wrZsB1xncWfGE9wql1vRRUJ9z++iGiPSQGxK6ogXBFmRP3jJO/
PyutV+X69YdVTw5KJBVCjp+Jk7IWryK7ZKXlo/tFpmo4ZrEjO4q+vFvdM4UzphPx
qYQ9ph7uvEByPSuYSZFHrOSQ4k6vqhTtLE2K8oZrsT/ZQakfDGJvZrMh7SLu50dM
1sqwS1+wGpbSUalwP5RXtQg1ymDUjAAxDf0qvTIWvJN5MwA7ZEZ/SnxfduPKLtWb
Y12v2zL7CxSNJkTuBJIhIE4qE8LPhTMPV9W6lP+M46yMsdUkgV++WwOVSQ2gINGE
SgxTl/dxVjF9b9tYHhun2CB0t1M4xhKK1F3X2pGs++hPW5Mk29AO2HwmWbO+HDtc
3SHW/jgKN1mUwVQ6Gxw6Q1NuEx/hKbOw/JjgBwMHsNr7w0IgxTXMkImSndxRecI8
nfkDWk1AZT8in6kIEuZviSD7csFdwRG695kUWUb5iWW9jGObHuXfHdbaJVmYRvH4
Cjk/T+SCpGI28wb6bWibtlswyBfFctPNUTjkRhbuAYLWzXaPyvy1i/FRjpmKnui0
6wtwNxoxJ2f/S1vlF32D922JmwI43RiwonANjNlPgtlCoGKqulmKQirO7tX8vWs2
r1czUtsLKkXXD9XAnV0iwiM1T9TU3O+6TQooELRAUQBOT/GNdbkNJdrTbiO1ykYB
zqC7lHiaxo64gfftmYCtAszrJt7YUD8bCDzIa+Nd3HfaCGoeab0A0URjClS9mzXO
1q29unHIeOCjy7Yd/zBQwpMeePbGXzMWKP8bdJccVwtXSJo5qCPBd6qnscz+Fona
ahJc+3lZXajT7FMn9TooabS+7wdhrL0Q/unyQEWZlLy6OctaAq/4DHKN4ZfwATsi
kwVgiMNOgyI+yFXecqmxzn+E0gfxOnLLpL6uJTwpMVCHYjV0L6G0TUULWZOs6mnO
VP5aoqDg/5oRDW0ug/fGDvd5B2G8PTQypQHbJpGXLZXxLQxJAYKMZP3BaBsB+Ohy
Dh6xn63nmlDU9m1dbbF6sOD0o8jZKC4gXScedA51Zo8bxO6EUmUczWgrwnOIqCes
mW/4L6TTttzEYrQE6WLO8pd5c267pPB97hjMtfOrysF6RutddFn9Em8nwUao62nN
NhZclExc5yJ7crPf51O8SiZpLI9BuQh+AUsiQNms8Gs7rDTLDY71qLjeXM6PqH2x
l5v8AzhVSCo2tQZas6YHCON03HQAgxDFZVgSOZJKml+bb6i/jOYgbz8ZglWBwgzR
n/YDA3aHJALO+riwIw05V24AeNGmSwgHhisqwZZqVmIbTcJNFuupRo1j22xTWkPz
2I5yQ6TQtoaZ2rn3cYiGglmnp+j+Z4Zwxcb6onov0GPpfLbOCtI/f6VN02Fkitor
WWOhaj4Wbb9gI3X/Fk8/fpFFPXoyZKbFM2nPRLLEnB1GWhBsWkghPqHt3BQAwQ7W
mLcRwv+jZvtRpo+He/a4wFttClhv9EIFimQdmns3pygDsQj6aTneVq4x6HHw8E8X
WD8ejNy7qA3ZaUHRZABd6I2hD04wKrkvpRcUuZXbTRIJWdM45SMpG8F5WwDoOziT
yUrVZcWyds0x5VmDO7hYXp6H2zzmbC3/NW5PS0sV9TMLV9SnmfRvDMr1Br7ZKl5Z
pHCMeKSqlwbLDkIoqQ3jcOawutiAqR063CTTuQ4gjQO13T4ToiU7K8r197evOOZv
I9fyKqnUgMq9q9kiVmWyt8/+aEGU6YWQvIyx3o2Yk5iQw9uuj555691CLz8ybriz
iGiglF2c91u2tGDJg6/A/XEXJa9dfVc1b4YvzYyHxaozNNiJRs4hIuAHjGArAv01
hvuvvw1b5aBHoyjEWZZHpeYXCRWmqX2nxMKnHwFuS5iTtvJRzgo96fsyM9zckzzH
ZYfnZmS3REYxemoHFHZkH3M/xzlqznO+L6F7sRX4SUXr2VdgXCMI/r8OnK3myzJh
JYbCbsI9Cb4SdNUTU1XYku+GUqzQO5eG0nM2GiW1LNAWe/8A1txGMeOzI6rPHU10
V1NLohJRzW6gd6ZfqE0Ok+2Lc6ohw+3QmfHKs+e5rLPfioO/K43JkGB6FBx/djAq
zb/x4Ft595oRcM3fCMRSD7RuDKfsSJJrS349xdBmsTWISnkRLYMrEQJGM14GH/VX
NLzIzwndBUMGbejWevbs771AjPh5Xg7djylUjMYHDKoNu6XSWxvnirv7ay0L75KC
3/fLKN/sCFQTp/OdVkLwuTIsPvUu1ioKWU22n8z4XKNSCmnyycsUWnpjGuG3YcF9
idMmOme+HFW2jvJWhvtcMDUgBegh8b6ZpRSdPA12hbq/coJVrWSx/Wq5yPcTHyCM
BcUzsQrqNNxd6xIQA1a13PYyVEZxI/QI/yx6p0PVZOFIxjSWwE4C9PvYA1WqYATc
4yUvaWwkSMm21T61hqYjx7OlLgKCML5MKKLsIw+7P/a/AtKf3ilrkld0Lpoim8wL
Qi7UFmgORFe+n6EXVxsUIRJLh7cknbiSmAXpDaUPzizWrKgFyHMQ4m3qxdQJPAXK
CtAMB5GV272UKnj4qAsiO68fnzGNzI6g+ds1/TUaipXW2bIBOfbHoH1hi56mjg7k
GQlm0vVqtDBm4tG/LLTDmtn8JevhHOguAUTFd6rXYi13fSn0iCHdPWZ439AXLOaY
Ty623oTMEbfT2EJEmSpk6tZa9S7inY6jd24/TjBCOAnc+KK7BTbOblTgVnyUZO0s
lSFJc2aLt5UOSHe7pnFmv4oGo/hQ6G2HdXi7EjiE3ngjJSoGBLQEbajlKn1V71di
XBQVUYv7q+lcyjNNQnLlgvTNI6nvzYO2pBSCCXCowZunQGNasp2B3gKb7cWFdDhx
UvrDbPuN21PcCAwwmaoxVgdfyMeBk+nNPG31qlmMoKj0zHUoAdGYzDADeOx/j1zZ
9Mou+zpfOs1u6iKlQB1QTbfaeWt5/ldZKZtDcML50+tTqqMKr7OeMCALJruRWVrP
pBSPcBgIc+iTSgEnVyfDXqlbVzY+5bIQxsqI3Gf30l5TSRtpub3/faIOqQg5MI8a
BPgvqd/Yy7CbhFG3SQspjHz+X+ryjMTUYWo17blnvgpiZwuVKmH/i/47+WEzfpak
lc9AWp+U7yS3uZfvzp+S7uDo8DVAh0OPJ0TlXVqG9P6vF9ASSfOAgORhdmY7dTAn
H1bNYlQnXYGShcXNwaVxaRjGsXzMEZAzK4LacKXVaXrG/4K1CjvPP+CiggeCZgte
8guluGuIiC4Jn7i1SOuSLn0ULhtqFhDAU/hQVwMSH/nKjKIflY5WMSPmLWp0yM5l
ZPbg7k2RaLf67V+HOerjMSXP+pycX0QbWAHkR9BvFTd9meWobIyGIgbINKm/yX+R
gsr3eXbD3jVEK8sYfuVcpFUQQ3SHXX8bmT+rSHgcATW86pLmt3mYQkidYsc+93qT
xNUt7Qd9jTSnp0MQ+Ffnuqn3+gS5TO+SQuGEh8RoAMA7Xin/FZh/0gf1Rm3qfh8r
IC226DqPqRyAHbUEPALDXtk5cEfPe5wwDXREuTT0Evh07a+VDTdFHMaizOB/jE6+
Xfj0ca5qsUFopUc3D+OMDdDHrY9tAHDnGujunmdSBuQRaJ+VJC/w6hg7oFChR2Qd
T/+fYcJSR8XLXa9UW9xj4qqP9o2ZNhz7uCgmWDSVmBugGkdoGs5TxYecXiEUGhmi
nTJVqiWffZeSdOiHz8fC5jz9H/MPMSuUZhm7/3XKAgYeCV2bUiMnoZlKOmS35YT/
9osy00s/4XpkRDcDvcqFgO7I4JseMKuGqoID5AZjT8mx7JzX17dIXgM0xCjrIdaN
1AGN/tCoz5YIwzBWj2bry1DBWPWwif7emtyAU4hP5b5dWk06cGUpZidleKQH+GHM
fjyp7KXyTUYFsE80H64ufGBmbDRjxMkjDVR4jOzowoN7aRbAfKkHy7u0KvolmAdW
UPGIfjBggTccD17mCs1ZwvxqCyyNxrNuMFt+9OBZxNiukFOvkZkJaATGw/Yx1sLj
9HR9jICITi7rrpimiNxa6F6ChO5VeMJNihoYufS32AE8Cdtb/k4dr3/M1ve5TB+A
sXAoN7PK/JYOa6ixjZbZWx0v++qKNlfBfAKsENQcC9zlnP5lPby2P4t5ZSR6kvGT
iETY1Oe6CbGuj314meRSeSINlbOC0FpPva/AZIr3KSJggfT4sXelHxGuQV/Ygdi5
h7/DNvB5qIfGcNdnblYB3PHq9OP2VpXRBn2RqvjEGTBmxpHOnh2gSC1k7g7P0c/1
55IanBVHrTpG3cc6yIsy79xTHVPgLK81pOi9XmHrPtQx1dduybhZF1IeaTaQk9Vl
/DQPzESHSvIYp0MnsPMF6k84ijUt7hlAQTtMttkXBEzUV6/0nihzlQ/nn89VbHVd
H3/PhDgmJLdrto4fz2ZZeuqhOF3/wDQD8EgXp7nFmp1D4W8nSdWEx8f/et4hbR1r
C7XvdHgE6Xm5msCh78A11opjkB+QkDWts2J8WYOpNpbXNHbJGbJTUzIQ047FoVXM
gSgx79LMevB9+I7RKKsgFytQx60Tf8YJFaf4lhXIhR4JIcbtXPIQSWLlx325oFS8
BJXRZIGwI2Ilvl/+x/GEjM9bgNClVDxJRZUcvrQgyb2WscOnCv4bHYCeETT8fLYd
HS2vKOI1GNloB9nbC8lhTBpFZEg4ZP2k+g6ehPqlPsYzK5ZAM2+Yapep5XtLwQNg
aZUBLsKe7vkBmehFxxavKbE7aCl568jJhcZ3/5ZwOCYXdEVHFoy5ic3cSIcQyrIT
s95Yw2pfeK3Q4kaHBDcHbhFvUunX8MnXxfAesT2zvjpZO03Rq3HfUV0yM3p8fp9m
O9Qaf1ydJki4K8gpCv4cMOhfCOSnD8bvQT/+S7joLaVdEUegtbh0ZUiF3P+Azsd3
768S8yYR82CNfZr+pibqJ6uZuvrkoJk5oeiGniQcLz1a0nuYXTxEP35FyikUHLxM
9mcH9nM1qwrnUa/r7ONO5XvDWFiZ3h4WuWFcjL3hO5lbjOfkQyXdfeHg8ncDcjAW
4l4vENDpgKJfskqmkjMxz5BBlbpPMI0XB1U2EB9vzgOkt6plvD2ca5rhjtYVQK8n
pt9zaF7ZfPdOaVyi2cOyWcjXfaqtb5aBpajzhC2wFrVzUrumw82zvEm194YGLIDn
muW7+iCLfyW3R10A0UIYyYU6tTgnSbm1x1Q92TZlogr3EH4K5oPyokRx5Z3DT/52
ViNT73/zZcOzvADsDwogWVFK46HioIeMbBLWVRnViEowwFYn+osKq5Ch45o6LKGK
8W6aBQVNegIKXu1gQokoLIbJym87G2/ZHqHzngMUmTLMjOvsy3bl5LHGl1+4Fe8K
DlJFBRFouE8Ns/0fsCx9ITxywjBnVhkxcP+4QnylsVZjBFgEIhaArTfBDDxpz600
uYDeJsx6qRUwXHyCBmFR9+00AlhmYo/etnD2R2OWAjDCKLlPBHn4rkZg4U7bfJM3
+c+NIuBC1OtreFJ14NjdTvcfLauVo/pMTetWszYYOmdkaGuyU8yRButkJrC3Zyif
rO1BJUvnpXEJLFZeu+VzTuUnk34KhK7ewD4pV862XJkW09zyDVKXRRJ1hG5d0cdw
bb43Fw1U/m1uBUYZc6aaWmn7mcZN2izm/ROydHMIM/n3EUEEr2kfBtcGbpS92FKX
kC3OXU14m69+dEqNa2FGNYPQyGuRXHEzPCl1TC7eoKBlInG42OYkOrnLSolRdxxB
XJgFzdCcw2t+/xCdX3X7AnqA9YxFXIRQsz8MHjdTrGN9vx2mz9Fb4vsvRZbBRcAI
zpNrAraSI4E2wl/6O3tZo14143nrxUV4fCGjnEgXz236wTBj/Y32HjlReBGP2e1I
hZmgz29OiZ2nPdexxidMLw10ZrwcOz6BZNSgp1QDo3Dv7qUiHbfpMILVvBKkziyL
BQkpvfgMRW4oBb23piuimc/yKkDvjKmzbCM4V65Erevk8fER4Ewmp3BiKMVYyjUR
018pRzZMwqpdiDzpEs4FoUyuNnf+xkbqUvI6qThe7u/BdIQtUD0n+Wa0OIot325+
VhLpiFNFrqlwFLH3ErOfmD6EKfNC2drbdaArSX2KUgd/YtNcaX09EMVOTm2xcP16
AWvCq+2utWAYGqVHBA7q4K1k3Qd79BlPxFcfmW7nKV3XcT5TjSJXN2pvnFzeCC0K
jvEE5olGimhyOcN3lM+8Js2UY3QNZT5MFuQtsZqsngSWPpgqc4Acory+7vTCsWFV
jp04y83qXnQqanVpXGzihmJh9WJuEPh7DLL1/PBVIVfQtKNqYxwcyw+Gqm/kEVSl
mkHzednEuSykMwIcng5LV+hGJLP9cyDwjDmom6gY7pQ2KwA5GFbfzMAvCtDXkhlV
PhOMwmq0D2aKdHke4VhwCvZ3VYSkF2sg36rl0AtrORsvETHWLsg9hfhXk7uGp3B8
97GmZ32nQaCssLMAodVvT+ST60QDYWE03iuT4Sl1fFSvkY+s2zGTNX+jnGagFqBm
9ZNU10fraPGrt3R8ybrufZ0HpFr+N52VcFLF5+Tmj2CKeUr0TX9KEHjrHhcj45SK
EE6jm1NkwyxlJMvASOMgQsQnXH2RGLNv2zu1LIpL7p9DqGiVdebmTFX61fGDreQB
mshnJJl6tmuGArjmblr63IL28+o44yS1kaX9AgSnVBAbP4+r9JgdXiM9JoaVrJ7R
ZSQdNDD5k3J/husYiWzsxALuyjaaRMqI49MG9loBMX/yZILEgDyMmwYwIrS8NuZT
X8adXUQB0MOatVrzRR7sVBPsPafHybGsGLQHlOO3ailLqr/0Zx6Tc1Tt0zdrlFXQ
as0vmQ4kiGCfKzNX/lndWk4zjVDjG79AKKyc4TryvOlj7656LoU/ud8fQAFBbxBc
AwoxfsDs7+QgsqWPRKXlg9bs9bzcCb1dDtcLmDgIAA/ko23y7CcoMMXqGRvvHmIt
mK5eWqDw1seZ3wZ4xA8XpW2sioAqdjVVT+kI3BNhjmUh2QAvnYJfVxYCwFP0ujwB
LksvoAH+GOLkJ/DIWfLWopXt6j+4+zofW2NP/kHmmRRyQ92CrII7qbhq2KIw6sP0
YersT2Qqm+uREPB/o3IS7D4Jfvqw37aZlDJDxQ0nfRIcVrTD+omHKL+g8pRl9kxc
I9G+8iMGbvJQKNdfiwSed6HPiuaHuyMs4N9TZy08PR3J7+hNdm8zgUazPcT4SJqV
cGnmr+8bJzr8OJrP0pBki3tdS9kE4z8ED95WelIWeNPMeqS92uDJoFkjHCNls2DT
UWEm5t6xWHUilGi9GEmW485a+kZXjyOS/0n33jtwbI8q1AZZdBMUXiVcZITdgLXr
gwccYuFRPtn5lyJsWOufVKjEkJIwHnidKn1I7VmMY3anik9UE4MXEneUFn3gJE+b
Yu6x3hUnl8KX4MVU9bR0r8oA6LHYZB/4NcE3YJJAbyXxmaT2NFfyNG3YeAu/fWFn
H5OKuGBLGuKieIDrT89ACcPJEhzZVBSAIVGhVN9Lf73dGP5k9+zAa/khV88VJ9BG
876t+Vq2ZKiwwZdl6s7AO7oy3EVFP8IXlEeOoeUySul/fOdNdBhtDimU7o5Jx88z
AFDD+G8K9cfSnG1RsiqnZ1c5y9lyYFlgDY+rfa4Zy6YpNGC+AXQKxceBgVGUBy8m
9JDgnqeWqfntVLTp4pN3NmYOxG/hkiv1KfU/kqn2mtw4OFGVB0cAbJ4Ozdvm4aoN
Rwv91n7q3DKI/QUr+EYp3QBQ95oZbWScCNVBIel68Pp8DTGxtiG95kLgqvTPMxX2
+qIXnZphuywoDAekpeYA/GjtV2ohgJ7BW1vqkCKBbdxGtSSZf2MlQYoXuoNDWTiU
+RuAJkuBqwkPFJQhfg/9msEweHe3J3YJQ7rshb/vGhM3lgJO20A/6lfJ+oNw57jL
ZBZEMO78OmX4tkatFWyWn2nxAVwk4w3Bq8ROGuxLgJwUTxCWxLQudS6h2IW2eRRx
DLOB4lUPC3SG0wj6hf2i7Ub5+J+ByC3gsLQZPrTtbaKIBJSUiFH9oDFExU20Gw8M
DLTRTFfRcHcD4rWMT/ZGUiPOdms9SHKJKNvTinxfw67g6lUq0H8tBQWEa9+bCqih
OnGXgZRa5cPplk8vpDUKz/sByRVl25jpKp+cJbmKuv6nmsTCYB33ssu20oSKyNS0
1VDRHH4OsN49hvwD2vlNEAcN5ZtEASxXIB62qdCPscILeb7OULZ1ypp331sGZh9e
JN2C4qWgTU2+0H2JInWt+7pqliFWur0kNsNJNzk1JJ5E5ANzSeQDodloONCVuzHL
RtTAT3rbykm4lJFk02Y8GxrBiQ4eGSD2ykbsFcIp5XPVX7cchYF+7XJAnkVMxRPv
pvNaK0x83P6Q8sJl0uz3gYQFg/Zs/Lr4lnJcFHNyNn/tH/Uq1HZZMDKMoZvOkYA8
cb+8y36cFFtbCjPFOPFPOdWUtw7JwD8vdPbdQ2zO8aCfxAWn0FqYmh38adsNywmt
tP/I5zO8GX1kYA0viaiyMvRBT5jWy37ZeYAgYV77aRJvojg8Lf0A0L1qs+jI13zy
fPjQvGi/fL8TRxjrb/GwlHXjjgzfmeB0AbMG/kkRpy72+RKQHfrq30exxPuke3qq
+OXJGHyfZz5c6SYgPVdbK4E9MSbgEGsrT8GleiAkhgqC8jQppmZt7zxP+T4MBn+A
ES6CeA+RI70V0cXBW0TpX3MB2cgLXplaHhz39l0939TiSX+wKaAPGdclS7FSDrs+
JTEuiKWGs5HQsuiRAJOHQ/VzbzSXcJ2ecJ61TmUqqF167L4vOEZNBNpUIsnTFwgA
WlM904Ag1b4mBxmmhJuQhPgch8jOhyyQm/LCgltOd1UaLwMTYr9wrCBltcfJZhWb
PjRHxNz8hAmilHp7iwI3bKToel6m8fN2gPet3PJ/zxoWNuvBYlpDUVPMd/hofC4Z
gMyNZ6+YqSV1EsMQcq7uaw6UHNHm8TX0ZYX0qaAlqsT7aI29xXcl64MPBqbKAESs
E9wCRfAUFkxWfwBlf6/44ahIyArMDwocHYWA0kDxv8+4zazxdGcBUD45muXsyo6L
7SipyLjmx/Yq3DV1+gM1Oa/j6mj30UohKFhFmjJKLxHFjXUSFrBXm2nmVDDUGwkZ
+yZbakL79ucERfDN/LjifCSUffYaHx9pY+vyTw272HMot/Be/wJ/Q088N+rJ09+5
+Hmz63RyJeS6cWorFFlW8swMvbgGXdAYhvIGL1yzhaSy2F6Trsl0a0tfCjywU5eF
ho44R4G1Hcdpo54Wd8BnUPFhvhX+HWNjuHhRioVmB7am2TiclLggrOpI1mcKzZDq
hrmdeGLdLOe+m8okkMe/lazVYAjcpT5gq2EtnPXui0Oize9gHVNvrEPEOSFXU52r
w8hxOXSs2qheL++YBL8QZkdbNrBrTlWlcvKDAXR1ZGh7YGip/ubh0iN9emCGV9vV
o0xKCbwykGEabwzghgGQk7Tvok7Br+YjVUGtVte8mVY+4YKUntH736J8QVz2u9l6
FyX3U/F5KD4nqYSD85E3ss3vwGk0ivkyIbtxIISpBnSpvzy8U212mDLkaTmRtwxJ
U98cw6oQCI3b8cjnxi0+2Q7H0zXfau8atja0HQuzU3qCXUrD2Yfyh6Tz1lssLXAy
P6wwryJgJEUsRv/rJZz01/G9D1uRayC0xWDLVm0DlhSMLMahyxRe7KkxDBxeijF+
i8fn4cye2VkUrlW6yZEy4aYoQhzMc0ocQSwrU1ukWj/bLSS2NwIougagkGJK5dS2
YLOaOWgWqAu5TGuFmOpPg0iQ1SHbsgsIeIokZ11G1oSKED1PcQL5YUutUc+xa8Yg
+TqCYN6fXseKehzPJQeofQdFO9Ea4jHHN7tqDSmRqcgZlCt22qjZv2d98VS70J8m
UD9lne/6Ofj6OAR5C/7Wmm6FLwKCAOj4wQTIoJv7/P5aAKmZPrDAvLKCddwtOdAw
ZdywEOi0WO5r3Qm3qbLK0fbntk9tSsxZcQ/L+vYtMLuQD8ZuJvj+obHbnScrA9Cz
EmnpYRLYG0uq8LlgfmPS0QPypkwgqbPvPwfDTnjrKiS5rTKGbmxVFcKIUVDPbBqe
j+l+MN4+4ZvYMdTLA/3tQElSf8qjKcm356dPDDSGeszFi+kxpbSC11KE0yxPZBL6
wlH4YK3NvsE2CBu7OZbgqtDumBKOIRlCzFJJCJoBzX4Ik4zioWQOv3VvWcPHjzSi
jrkJnVjvRYZZTLfDcE91dEURse5RvoPxLp4Gl1BV2Jzk6o6Pq7eg/CSoWtK2n0Xb
KR3nanvLCrCk5ijcaB/c23geFKnF0eN67LS00Fv4D6sz1bbCE5BOlxIPUSSNqW3g
QM8UTiJ3GaeGaYjh5jFWGEi8pDBt6bN7R6dvnGhjovUB+d1Bh1M/VVZSSw8ZEOqG
TVQKejwjVch+2aYxAPYNVJxAcz+CQJC6yTCAa9ETcZAPFhXZQp6DKXAftwJkx5S0
tOE5fD1jFqfqr+Ajkl51XrjM+bXOWJk5Kers42oaYaENNOHpjtE6Cl5IXDAnG/yr
9dzwlL0iDCQqoqZl68FQIrvgbs7P4oVUVI9ENHCDuqNE/R5T/wfVwf4zlcq6SvL3
S2GYTC/NJOoUcZTpdAho7eCJOh3jpVos8hXJ6G0rYOZ17VLnGk9FFw4zSzPCN3U3
ZTYr2kXGi+R7PZhUrgeQLF2R5XS1bssqabygJ8P1YyJGteEfVhJyKV5+oQ9ERYrj
HPG3c8AH3UW9NUZO+vhtAv8fWkuWUJPfwpqIubCdze9Iz7YPcoHV2MBcRV4l1MzY
h93rxaI6BHiPVsInP3UvhsTkVhiRFJcJWa6xLOyyYx7hWW0Dkn5OCLDyjY49pkc6
o54D1X3iVzaH67ElV2KXGtslyXEOFor72sPNcZktUKPKAbtbFZOtkYYzTZDPON86
MgdkQAjw0wNUGoTNVV2LTayZ7f5ZpIly83Zh/wl9ohT7u+UZzP07zEO/fNCwgc0k
bOGA+0iL0tthw987ic69PLhRJmIMfYTKIlZhr3e/eqj0MdH3VWMJmc+W+kfK3IY4
NPzXWa13u20QC9XOfwqPDJB4a8e06Yvrgew5EKu/sVZfFJilHyEBH20Jmr513lXJ
PCnpL1l9a4qcznydB3fmQg0SaE1N8xiIU1YD43W958uUPSRorjkFOjzl51GUW5zz
BJTM0OWFQNwdTV1J+83TjUzc6owDrBX8mndITxRAgG5ug48u2kgeBxZbrdI0vooH
p3/kexqwRboEm/p4UeqkMs+u+vNysCVnqRFldnwmf0Emos9FDmBXqdujLoghhbOD
jfE50cl3o69UYkjmurZvsuUal5K//rwJSHUPr9V26eKShK3s+cfzBSA5pnsfaLLl
/CkSYoK5L4BAyNq5HIc5DZ8vEbenQfIcu0citX57i8iS0bg7TR4oCK9IraIGR3ms
BibyNBTsuObP6lHtJKjyfMII70da+eCi9mZntrQCTVHHa5dEDXvKvgg/B+riHslM
uORIRhJj96N/zlDd+WiPAWlUXwaVL4fdt9BKQ77u++9z6QG62g7+nlIrhDfNHP47
j+K2NSa1YX+Z8DUt7eYMe2ITRfgjgz7AdK1bJ/E5kBB/jiUtKdyfOA29Aycj1J7e
n9juDyxbMBtbKly1dPGlEST+MJxLtLLPqVkmA1Dsq2mItkpu3u4Vu8/q6YKlDugX
4DKqyb+94SOWboS84hzLaUB9Ce0muOm7PsDg/0IiOdn2kPlcujzzQMuDhJDks9Ac
jtAqrOJIJJWbUoxncTs9/eV3wgJl0p0xrpHaz7IzRP4uLadFAxPNjHabglUHTeLE
2oFjEo9jjmgw4L7scfF895fkYKGZboRPTaHhstORpmdu8WeQbmTJpnxSiJrkqqNb
UakFA8dRoNK1kduX9Q4Q7FZG19g5GRmyii4CAKuoSjUa1+eH/HcuRk+XycNV8tZD
jqNXSi5xs/mB5D0blIXRl4weprbaGdJ3+t+I+FYVvAcKEsLm4wKpoSu3t4NL+uKa
91Q5VPOZfX03pkB0FkD1XTCBmAGLbnfqvqzAEi6cyKuk3ZzOFMk6UDdQomOEXwPe
6FUXAMwCPhxGVitdMcCMXhgBe3kTtt5AfOmaPoipaqTFuAnbJc54VLhUCeiiux5Q
WGjOUdEnuMwVM5iC3wHYa3YWz8wivlA5EK6RfeNsNqX6NgjGJINrk4BWGTwBWUDe
IZqAw0nZEY8TunBYDIteTnirqdbs1dhSP2J+HJbQHQNoqXtkfr3wRUAzhONlTc6z
oEWerUgoTlxuzf4o+7G2qjqH4ABYMpb/+rvnU6tq+ezzprEDiYEZSBYCqrVlmsV5
GfPuavHX+yPxxYa+da9mJoPuFsqmUmNu6CPWJjABjVRKXTYGDhpazyd0p/IF/wMR
FTT9L/BXgwyVYEXMk967+qECgxX8WScx946hDHt167wBrVzMZ3JVyceA+weiZMZs
xZudFio0JsD20urV17HUvsYP1rEmiv5UcNrqhabfOprfr+DP4RgNGDgRfyqpWL5V
WZVKq5RRCtlf3jvNSD4PlW14MfptzIC2t73ozrUVId3m1UKa53fCQBrybuJKwesH
5jhbTxrpMTkVJ/EPCc74XzqWCa31yDQmS6tRVcs7T29qsvflYKPaz69VSICJoh6w
ubrlju67HDvl5fFR7TG/CMDUoOvGVvOxRAt1UihdRZSlTncxtyT5Pt2L5FfY9KvX
F9DlIo4OpZZuEnpzOUXJGz8fcdROYc7qQN07qJm6V9C4JeSxwunL5H3puBDzyeRI
0VO6EPsLy3cn6vxKM4TOLfVCwEw8Rj8X7Ornt6YoreSUbTKcveQw4LXqF9G2yZuI
3LD2O0i18FCrd4piMxeJFlw/lzLkbeZaZKHbqjsEwPIg0X/AON987MMiF7L+3ZVv
nO33hywGq9w9cZHbudK19z2jzYHFa0uhEW/XMl3gXQh2c+unUugciI2KQAN3zNO9
wyh4493Fy5br+2fPC930QPPK0ny7nhB3P1ciVKxCxMJifBxT3T6hYa/g77xwtMl0
WS3OaBvbGMKjY7fmYjJiC/QDm3bW509PpBbg0RcZF17D99ArnqOPisCtCTALXwxl
WCtI4gzcut4OolCsAeZLRvsnGOjWOR9v/ETzqJ/RZgIqR/qridoImnSUWvZhuxiY
4dRD4CDu9N5c1eH+mFY8DAKSsVnNyX/SECOMCKSvjaBpATBrufZ53VHkA/ck719K
FOOsLI7ogMRuKi6JqxG/x3mmtQnsf+HQXOevsHCclExnTW3JpWq5fYi8TPsUUoUF
5uRqWTP2VnXyovpVtm+luPPMCdu107hwyT6CZbUaF1pjPRvWpa5i+8Mhg4jCOgtu
K3AAfFZUqZZPWXQ4W8Q2M1Tm7pTB43WyJrDeHf8g04nqHOkHmrwRWx4k9KeX6aUm
uDBGKZ4tYvrhYHbiiZIvO2SRhkHiKH/Dwn189x6JMl+sm2zXYdcb0mKL/MkGZTO+
v5HHwTKi4P3qd3+3Xpt5Sm/iA4nvldXj/HYx2RX7tV5lk4uH6lCOI8sFqaXkIP8M
56uleHBcRotyra4nL4zEWasgeXgsoHxIE/+0JKwTbiybIJz4MmvZ9UUsjCnnljZs
mAlq1d2VUxdeOtW+KXl0WYl7+v+dQIr/ht/fRu2GcwyH9QgVI4OtsAPlmAj/X2HR
JkMSgg4lYhWP9KKN99AMkkIi0s2P2i5wroz4JpYm9GFl8jh9VmkERaEenJeo5wGu
mdcCJ9w+WXfJGYL7/LN9BymI8ckfUsWpSnbm0VOzVzxFRWVNDQlPPdq17dojTJTe
dzWntmERp/bjjO/4JRJch76Br/kaB8eN+OrkG1lWtAiS3j3K5K8hHeans8UPY8AK
KeATe1cdnZFcvvr7+ayTIN9I26KRGt65tWCYJuQZ2FRAUk+tgYwqFmkw8WmEZtYz
tjt1LrrxpsnIUUdWEdXua68BVOiG4xUy0bDkhMiiNOsn7484F7Wsg1JD0q8XLtdt
4QA5qIj+zrA/o4aQNCHJePWILt34Bj9Wgr0safXHbs+VtN8H5dwuYt6v29GZpmn0
qZJQXx49ILtbwxhiNaZjIxxqBzoYBUlG00G76qheIYaNi4t92k2O+LwQdgsycAeJ
GywNSxCHlFbCE3zTuFWyIEYm4oFrlfVdxPKvxrmu9MYtvogPtIzW0sAUv7srJff0
Dhlj21FO26zpOaIY/Z70bb+85oNXqtJHe2Rub34JDvY2aMcdIRNL9ac4gKg7FAS1
ilaHZoL9znBg5oQAJG2AhMrD1SF3chVYW62NcGj6oFzyB0F2rUltIIE8EmnaA+Uq
NhgQnxxohVLzggkQk2UC0OTi9IUViWfbVPCyZm0pu+uJ82QrlECCqL7DGIonLtah
J8liRRBx9F0f3d7c3wTNpbya/Payg2caYD9WtiBDUeKEZVNUMuJk+Mlve9ninls6
ZOdaAbJ4ny8XV70uiYTFCKbkH6oyGktu7eBh3zfdc4etDsEnA9yJJk5eel/ai74m
jCOEzxNNObLqZsU2zUCrvDydFBGW4UTmos9ySquIBRrC3yYvX4ymfvjuewvfn6tc
6QTlsdBrAm6e8NoWLU+PDqju0hesWG6xETd7rkznQq5P7Sdzxy3tfShxroLk/uag
f6Tnlb0kb1AZQVZ0loubRcJ0Pe4+SabozeantuE/IrP4k3RRXMD7AIbjorGESjjm
S9xeitxXrWyE+QRzL/wt+bnLDnmQ+Wy0ObyG8tuDuiFrOJaCBBCKA1WkfoV0aiph
tnQoqQ5T3PD4R3x6rorglXDpXoGoZsfUBR6vR/og1+XlbttnB9PKvuamVCqVcnEo
tQ1nBLLc1a/m1leRj38E11SuVJi4ikHYDELi8PKgN1C34QP/A+OEOGRt037TtJhj
W+ToxRGcc+i9ipru1eEtNMcwL6bQIivo1ooMlfYiXO96LSD17M4wzDRQE+zVNrMm
cK+IiB6xLCk6Cjno+fBhcxxyDcVpNLh5edjMnA97YdF6Du3sijU6s65zFbq3PjYB
NwlJV13ITlLabuhxZ2vYlHvPeLzf8Xv3+0BTtPow8xh2Bt01SE2gv1Q9TjAWqV7s
766HfYXmPRmMoSLLhlbjfzr+o4k2rcctpJTIBKr5Zq63D6ZQCnm3/MglKOpc/s3F
DLYdpOuGvUIn99yQWL3e/tcq87lCpPpitfTPrJiLTs5lw7Y8YGvlI0rAri2zE7nh
Ty/XiWlbHDpgVAoxParxaX+18RuGG7M4qSQ0XqRwF1oyvukaFTbUqqJS6BiVGIig
uqwHJrVkB63r5cTBf4vVn58muxG8sf42t7C4OUT93SL91XbFYrDitl8HDosFgdDs
F6DDEbbs3v20lgbxnZmTUZTJIrKvSyvloJtqhkmctrJz30naF7gfeWJMYJkL2W2x
I1KJ+yFY/7hTrPbayY0L4NYPAeWWc0CaXkgXdXdd2h3dLqiSnGMD4DAB5OOg3IX4
j/GYeGbGxx7ZwEucYvYt/b9OKrGMpkdZDcsuUlRU02E9F7/+87GE5T8A9BP17A/g
wdfeA8JEgdBGhXIUYxd1BTHn8cxYBwlFKOfP8Wqtf72AYsHh2mErKamIhr478vy+
EKL52jMP2fhBtNAfmVE2LkUxdI6YVr5gavKpuk2pl/7lcWNnKfaEybq641dAvKqS
QoPNg3lSKqvG58rwYd3CAOGE02zAi40uTptDgHs03Mr48Vn4i7YjuvDl+sqqVK1+
1AQvXVdOzbnjwgvxNveZaocv5hR93wSNA2qPW/w2dY9/c5EHtj08omljfuXhpk3P
SmldFYcYHpFyC9lG/JFxj/mrYPboO6BSD11TCmWooMsussAsjsFqjKhgxsrpjELY
TBVutC7VmltFPVQDV+UNVgYv7b+ySgkeNhhrHHNJSm3n+Y5n3URZ5jLYnEnZNwcn
AGH6HRHl2CGFgo84GdfEKAHvGRCBcNrM7IbMXrv8cfMylJpYWshem654BHZhUn0i
GtLeDeJBFJrnpPj6tYHmPtoH85NK4LZlxGT/2fB/SkairPzIQPYWuqWyYP/DcaUG
8lpto7ydfvnLZDRwSnMWCebn+Hw/m/zdbPohmn0rLIHxefubBNdc1b+BgVERQ+sc
buj0a/g6xwsiAGEvgRWR9xEbaLmRm4sBnIcUcPC34KPXFi9vmLWnx6Y91mG1uIzI
9bLK1RqBi7mHgchAHIrkfNHGVP4IrQm+MvRo+vkR/sKgd7LUX63z9FxHOcOz/p5S
4HAvMSIxyd53K9D3qL4HXsozI5tpc5knGwgeV8gJYaM4QxrrnxFr6u/b96XcK+us
OIT2FPYuz5Uip9r7w0Dp+HHdufnwW0ZjzZi7y2BP6bYLsONYxUTQYj1nEOoQVNXN
EQx8DRZl5sbUOu81yBM4oDuX6BbiMe1Q+Luj7nYTi9QEkXziUXxcrC6QSdCSG1q6
6k4xRdWXIIC6Z5+lkyfGcKu7EE3GhEwHmhgQEL99lzq+yJIljQa2oFxP3IjfZ9kD
6quQCwECO05uGyahJggI5nhGnBxPWDcjRspsiNDn/IRPSlpl1pSS1ZusBKCKlOdG
P0Iij/ElA1kB0AcN9PQWIFOC9IfTyiYUTvBsdZk5Sg5+07XpIvpEuwfzQuWflWfs
ypGCULGRRwzBfTTghd/sRTPCBGnwyZ2CQOJBP0XqA4xN08eeWHwZzqyHutv+cIpw
r669wjIbfN/3jFWQynbemB06j5WujZ3RNBaBMQ8x6IQvs6H9clGqsoHYcsDjdIPb
QBn4nTT000a6WSSG/e5tQNQVnTHkdbru/wPWXzufKngSxlZMUo7kTNQBarnjKpIS
CCqEAmN+pTxONcUYwV9LqTkafURGp0jCrUWaEZ4aq38HP3oydOHHHwZm/yfwjBfL
Va6sewlrwrkL58cSRy9AkccEGGiUuLuzQdFHMz48pcPLIrBeiUhFE1ko8E8uwUpD
/C4Yox3YnPqSSjjtBzwrVNx9ZadhKIJEa1HpNrgV3UidFcVkD2MmwffebkauHop1
XYvjGsrkInFh1IA2EOCUqHWfcrRXIMtU0aQQ+SXAe+tk1KjFdXmLFVKPl2FOcb2Y
qTIiJChGxjeLpPu2+mJZXdU41dDPEhX+i060hz277KqgeYMr3xFGeO4LUf3uOnZa
pmo0BODzy4DFf9TdZnK4jFbqH9SN0YQGORYh/FEtEv6IX2NAg9GYQRFrXYyj69M7
I0bP2gaMH0dJdVSC0sTR0OTYfUwIsYoVz328mbfvppg0snAYOR0dsxK2/5IHEswG
d4nxzh+7LNw6m3IwYgNsbROxEEjezhZ+Bohm7AeUj3a7CAqCIrx2N/ciQUcEhnfU
tp85+G6nGbtXZ8Hb7KkhM+8hux3GI92izLjz3nRxtdfh3sYD/cVQZ9e6jSGIw+Ef
ZgBLRDbScuDDRUvrNGeBE25MXSDlqadaUJ5AjG2+wLlClUkRpPq3a3pFfZdptzhp
URUwvx93Dmki8t9MdRyenUH0mz3McKFvNOrebqCtNWYtxQb3olihlA78wua+WZrs
RLyiu8ldISbn9oo0/p6NyKOmkDsNnHahr+RNDxbfDrttl4CV8/VMDxmes9/O9p/k
QsAFRcRgTf5jTABlv//dcewCutgCGAlFw47WH4DopZZkYb9EfuB7Wee+VKwE7xkh
UoQpGVbqGHFSCmOtC29FS8n90klyGXlPXgthReIyg53NNnPJX9O+Gl8uhasmCcSd
G2BZjv7TuLPPdNL25oincRfTaWgpREygwdhAy/OCEjIEpBu2dCsQJ75SlR2pPcsQ
G4Pc7cF1keyu4+05vKbXcj1g3UMF0SHPfg8lddVhGRUIUClmq6SmYM3oX7f19hDZ
E3bi8X15FqLdYv04KcDH3XLz2zvfOqzdqFWrryng+IOtOxAL1DMvykp7P6S4112r
O57vWz9m3czswsRu+ZtwzRslqb19U/06B88zc9eeUsQEI5x6ECqlBBGW4plsELnv
Yho9/g8mXHHasZdfts5nduW3CaP+J/jnSrlSvjtV1RvK5AgQ79VRjIP9loL/sdK0
JTblTACFZQGqkCS9XvUDp045TTJIl2LTsl7HBVMCjLIEGH/6KekZE0LFzlP9nlVu
xW1yyuuUuvQV2HGu/5P7M2h5A7ZCQsk+YZXWHVYDgdpfmDQyLeTbZn89+IhTiIAm
YJfmndx8G+eZGJlDltJRxfhPDdvzlVYjEe/OsVLtvXnmvRHqtvA9iwhXc/n9WQMM
lAaodhFtX4ul5ZQkZBDUEESCp4kctwgcgPuDWRcnTFdqTDRBOEt43I+YsxCaNWRV
F6X2pv2KgWFSUkOsa7tIOBgeTBfQPOUbu9Bc4B7kP2iLZ9OPIwMobvkFr4wySKNG
tIABxKNMSeG83yqn3C3lfyVYboUiCJjceK9iKdruN2eKNY4HSKuvuvfS1Sdzz29N
tXl8ryiATW2R+CfqENZs/5f1+h7eWZIfQBZ4JUuSMmN5MXgYVPGlAZpXbTsdiRam
Rla/DbEDWwNJ+aqJj9fHxXu/AtV8kBz94QKKT0o9w8kbDycFtmzVS40sWNq75aQy
IM+/ujynPZ/bpTCut94T8A1SIPFU8BSNUW+0vgGkSPJn0OeZRKvbjgL+gRR6UmAV
5HnG9mLKM4GZXr3fCCSrNRd1D21P1C3z6VZG2eo9xjqHQs4wwZd2wB+rl2yXTM22
32abB1AeqAx5UfeGRHR8NAh477U2rPZE9NCQbpd46B+i65AL22XDpYshUp0XATpG
RaND1K5VcHA+3xFifUjTRNY97ng5fr/M370cnDSQEsBXnULoBnkv9sXG4ggj11c4
tt2E7AZk0Ignq76eKYopLQQz9MzzxP97dMrx4B04XnrCBYjjQUu6NzpKlWR9gPcN
UFrFdVNyluiuqk+k4bz0cNhirRm7DIDU87pYRtic24S52Y4FLyCjja60aMvPhCtk
x5z1OKqaDHYilP0rYHm8ujMECY8zbnLVDvRCC0Gc3AmNIuOZnHFnomCOw32EySdd
mqXvGBVaWAC+XEej/RLm0sU3ZgiUREIoZZrdXe9xbdsvprFIyfO2f41yzxGlKN7E
vGyYQS9Q+D+7fkg1wDArt+dj6jpDB0RFIRjZD1+5bAL0NpW4N7cK7EASVXUBJL9E
c7Lbglo7o2d6kZKbKG09CaYyVCaqJzGTtSoEGz3XLJ8YvVMWplzFWrWw5WUJGEgN
OOmSvhQzjUi11Hj0+0RGKUFpTNB5jtQTo+mFBREDt5qH3tmImEMCaef9Nh5qsRqp
oWz8QvReqfKxZZqmNujPlfp5WM1eP76lZswidG7UV0R9N9dmMUglcMmWaM1cXjB6
bGFLuvBlWQWEXMX80DOtCFGNbbD47HWvKKe96iqlz92cAviqOkebP6Pat+4JLOS2
HGYZv3bTKOCxiI49dZX1wUTSwtnBhiuL6HyAHBYm3sNFrQcJmJKu47aQ7uDLaj/X
7JgF6KnxuZgTFLX5RF5ZLZLV5nOvFE/EHiWFkkqJk2KvbKUgIbrsjR62IJhkkQpq
mY7QHyjSzfLEjHE9tseq5lesicOA/Ha8YOq+xiQ2AzZMUGawft39vGzH5O+M8UQD
Lx1uAj0lULl3jOKllFzpc+l8VKnU/PTPMIJVpvbt+Ux8wlXXJlegq+HBn2SgfCmO
XhHv4roosNArn0b+7zwDDDpNHAZVY40S7rOKV+vkaaodSEsX4VNX3onQ8G4PjhuL
lkC3/JsKd57bYASvwdp/Wkz+iJE7LoDDi43eji0X1cJNrUfjzV79thon80O55YY3
F8RkscJdVREvK/7/L2kTqSHi2PJIs9v4SDg+vh2jdMGWnACILDTFl4bkvdFbQC4s
PKqKGCzBA0jcia+Mib+N02Ba4/wgh+4hQrqLUa70RP0IbUkQhbwybiKU7hWcG7X5
hKAa9yzO0EJ3BFV8DG/ZaIgsAavG7bobnSr8uKih/ebTt/sn4qSf7oTc80krdotr
qmDhYZ23SNnPaFKXx1985SONq+3EZf5RLp62DthlY47EFz0hO+Q3Ft+8tfpQNsVG
TOLm42bgf0vJWt/PpCcYLc1HUyqnZOPq02DKSF7B1HDgDnw2/Q4Q3pTtCpwB3Bd4
TcHxU3urAWZMgOsbTXm+A8KWv+UmiITVZW+8+3IPgPM2Yx2y3Nj4eRdjrwVmhmQE
usEBrCmMEYuf2StKyUpCaEUfPuq+EONa+EV8P2xYjdYuwxNGwX8bBMZl9aMC2VKo
JuX8EhrGU89ymwjZaoNYGwGlqqsg4Xbe6lB9CI5VTWdz5cujYmxS6Kw2TEdcsuug
O7G+bXsGuwKx90hIkomxLd1+EkyIjgT58DZ118PJeVM3domGuLARUpbBIau/u0jT
XwnCjKohoh9173L2MuCwT6bireSX4yBNcCbRuJ6RKcp26r2PTZJp2bxG4Sgrd6RG
53z0USZf5IhZyuG8XaGhBO/JZnKPmrCJ4a9RITnepX2aG6vTmyYZT9hPsyJSsNq0
+Ozc1qrkruEm7z8CFwJ0Hh+oncxEC5D8EXOLxZih7IL8i+zPkEOv4dmxBXi6+NXt
9HNnSFopN3HAMZe3NNvvzTt/VuiZp9jk6jsbIDhjDsCJmhKWCO1rS8/EeD4CFr+0
HEIj+l0QXyfn5Sgg0Ulg7QqyDwRvvQMEUWSB8xBsFy8E0he0jh0ESlruu7ucY38s
AaZ08kLXXoRMKHmTf7woB7MZYziCiMYI87URJ4WdqW/amhvE6OrBhFoCVn0/1YgW
HJG4GxFpZFE52W6HGqbwoJPlzImqWSBoqtKNHLUkfeRczJNdX3orFYJWU/f+2NI6
TD8CHMWmviFmHAJNT6L1iY5bEKmmd3DmvWCylfRzP7Ur8WJTFytujEG9zWMVvwU+
2CFdDOZKAGLVo1gSL6x+9zzscm4OXUg87yOqvggllfq9VZ4mSDrCtmc1MStjqHLM
I9YSaVwM9NW5nmwHqaVzkvUw+l+tPsOucjCgY2msdx12bETxPT0YSq4ByMC2448f
kk+Gj8rHSBDQOenRhj4qiyX0DRvBaJtmgYSrEXKcUIJvzTBb4446MMYiJFnsaHzT
ASkokmCa9Gh88X8hquXxKRqGVNVaCY1tT1HacC9mqDoUqcLT0bFLejFA/wmjR3vB
Si4XJ9L8LvUOhL+D9kCzHP3Y89pEnd6ng8OSAsAhq8HGy/rPa7roijlquYlhkQOn
dJBtTBjAuaia2/VD5P32zzY1s4uyk9QNfsCzzkVI4qnWSrmgDkZr7hxhd9o1junN
7DjxG18jAtrFMbGMnRR+uhF5ZC8igWnQIvc+5kDkdwdTXvOvFoD88jTl0Tt4DpjX
6vABaadS3PSPYTgRcga56eZ+FPRTwOFFLs3XVdJknwcbzIxWXeD8eA/KztVZy2Jd
5Svh3AaA12spRgef5ZCHHqXIAqUDk1mTGiO1zdwfHDwjhObqS67QE2+D3QWRMZUL
jOqBizb/oAIsws04cwuqwD19qxY//oR6QlNtHw5db5HvE74ao2ny1f4MkikiLDpk
SkaEJM5/xdWm8iLojXKJ9PneKP8KsIHdS2chwNyRWxziJAgrm92XXxogp41BU38m
OqbMEd8AgODUFfsP0l8dpW3enL+qHAnKXAZV86IG/p9UC+tl3LlmungiYgFFRAyr
vWr4H3MnTPl8CEN/KPf2cbIF2zvrPg1CWN1pvvjyCjN4L5mjgxskovp/KEfxueSU
lV5jyTzN+BEkcCk9H7pTokpmp87EC5TDbLhHM4MFvbZ6UCiIFOs0d+hcleWurE8A
1Xs5fOi+qn3jOOHpl159wkCUf6mf0uRfli/7iCnyatBcUMCLlrAcanXLr2dAdokb
R4GRNg6OLUOesUGtE4SrD8Nsbwc0SRaDtZre05AjeyenP1JUdKgqWs12iCetnhuV
ULwCK5OnVcgJs2qE/SglYStDG1/EUs0Ekr4d/RH89uesBBKRw9rERVog6vrNajnm
BIRjyVJHYGzzorm1dJMCmYIS1JaPftL3foWbk+hf1qRnta/1ER9BK/gifOjR8g/Y
V9CKe4T8KPLewSqgddV6LCKZ6uwEm4DsLlszTAW/OI7NtnAsjtAfagwJCVPYzty+
3fnX63WAAQ/BDJOsJpt0UZlDkFRDiHM3tlaMZjaO7LMvDdIYnE2tmlYl4fQQOPyJ
jSbI97ziqLiP29g9njrf4SMeXcrp/fjJ/qr18dNb03CkjA5e1fzQrjNLM0Tly2i6
tKu+jNv5AC6iue2+kWiJANmoDNgWZkuRwQMHwvJVeNf8Lx0qrbvBYRLerSQzIwSg
vZvGaZiT6/2TrD3V4HBsmQJHA0Rhih6c86TexBJy7lPqY2ccWBza1kzAdf0Q3nDj
jBDfLGqUwLaaztGlxT+RpsI9p7hh62YKsKbJNdQUCo3OJg0R6MmArxxQBVFv4e8P
9K3pBBD8iNfSymsh/q+F7a7znxBYFRC0DAjUN9sde5pGIInl5p7GyuytLpbGsH7G
quyVcd/rpqQJQuoXVQpHNoMU1FcLFvQvEBWoAid1kuM7thkF93PvgUabbj0dsRJC
uoZgk3PrlG2JZS67uBwTa89kYiDHOqHFIS6Nz19hsyHgiw4zPN5zZ5I3NZ9fW7Bu
dZ2ld6qjlqaiCWML3eLEu6VmyyksuRKHzyQL4YFCmwZvIOMzWcsVWy8ql4Ldoial
nC8+g8Ks2rtj2JxhrgmKZFVoJZ/1WYSSqiy+xC3vSKgQgSnl9SbKQorCwvalCsAL
tyKEe0nYO3OLnl4nG4nvTbP1M3S9R+JYrOnGYXEMXUxV8q/yV3rhEIsmi4LKzZh9
FBtQbr/IJjCLdadyq++Lev7+0C6g2lblCGGhCMfkgilbiB+mgIp4iuPa8EPqXGHX
wF2i5GI+ebOSEMCf7ctterBqrDFU6Xt2KOnSjZA2wSjiCu1RS7hi1e+W4pPq2hg6
1/m9ehR91XGCQaRLkuKSrd6/Dt1IdgrXY/5Kkpgtv1NDmHaqmKm0tzWNAtZDx5W4
1i6PYQ481M8IHApK8pybW5wgPvjIZfVlrbmf8omU3aXggRHzqck2bb5hnvBUOSY7
PvBPuigit+wFj/+4BVVb46SveTu1+LTdrE4U6yqKlLwq/XOhCAi7vfWEyBdNAbuO
72FTqMXQz5rTCToa90W8Q7SacPPcZxeKAn8PKBSR/YFpU+Gg4MeM6wdaInL9p6hX
/j2wWAy6X1DAYT1AclXwJDKQlSqfcZempHrwvLA0rdgHBnHXakj6kE2TA2YxqsUB
QUwN2gFpU0H7L7z5zpjHqWBbmULFUD4aL9l/fsijKPlRalJ4H/+SsSiE+j3BsyTn
gHVUjZFptIpeWVJUWjeNXy5ja+rYI8WFSit8XuHq+1kkzc0DrfFRom/savR3/nbd
A3pixAcPgoZCHFPfs90LTEpm8su9nOSX4WJaCgmFJy8DAtYWgvv7d+yc4RA+4ujl
EpcO6glUH/H2vp8X23DO5rth1aaYN+W0RbSnHaJ/KXZNtqOW1NGMqokmDcjHTOmq
Nnyn7c/DWcaW+K728d3vNCAXugeT2meGhA7Wn/oFkjxhZQXrbNNvjJDtT9tg/ZDp
tObBXLRJoCTc8tbl2r2uJCKCXm2PCGkupAlna//iJrZ8MGLOVtxscxDytBlGOWhx
a9k7zxi1LurRI35EiZfuzsfNyyOn47QKAKgr21unGN/PNhBtBgmJkZvV020yPg/+
fm22BTTthzfVB2nVpQdCb8p/iyffUck1bBI22td9B5TwGkdZak+ZKQtz9Lkzb5Dh
rUJEw+CGrHClyl4OKNYqU7vuS9XuPGzFya4/8pSRzta5hpihq2tVxYkwsiTTK4vx
Vc2E+2BtB63PgwW3JUrXorrtW6v7p4c7992Dracpr9SxtEL6WISb3UCY9D87Ce6I
Ob9BVqTf2UMl+EBm5J7PLzuTxvtDWhvd7nyGlWE4ZvrKG30m4B0Cr3H7B7sTfpB3
VTnLAhfJdd44p/4Wvww9/XoiQdbo1IFXGPU5yM4vrAluXQytcoZTLgWST0XIrneg
PogyhC1vqX7lBxWbuR/jp9DwFPfUhqyVBX2c5fv+QkVH6P5+PmGgin58gtf3f+wn
BOHHs6OWzCaCplx9/9RCPIFE984tNkdyTL8xvyODmWpJ8+cXNn8dFhGrE8zGmATz
SHyx38Mbr4fqP3lLWFtjX2v0VpzduZ/Gr2J0nO1XwZPe8eq093gHpWvqFlM+jNJB
FnML6lYmuSIZK+slvcjQkyF4XFtuln3AtqzVDX9z6bihRRg1cWz4eEV0n4s857qx
5xLldaWo6MiAFHCHiOIqg8AZrlCEPMdx1hnjUKnFVvFRiVGmJCf1h1P9+EITnc5p
I0Wg4xn86Sg5m3Z3VqLFvcv6nh2jUiRuvDbPd78LqLh2w+atBrAB5VmFcqoug2/o
Af1FwQmAXZTJjWInC2AZiSEALpT6l+QTAHBGu4WmFpBb7iCm6CQywzqbvdx30Mgi
a7S2Z6Qqz01M7aWAK2OcP3I7KBKWzX8VyoXvo4vbLlRIFYzlgc/ehVoxSXDkxppI
fTFvWx+fkk4GPmPZVJL99cmckZ9Tko6tlWePvLU8WzaC8gl3xB6ZmigdeCL3FWxP
ZkmlCMdSNGT6v1kmLTHROpWODXcF0KHfdW9aW5qrhWw2r80ouCqCMpKNDb/FERpw
SSKrGOF9/AITPb2rKHVKwurqqNvzH/+T+ScUiinUpD6QMxQy3h3gjmw11WZzmyju
/ubyih/AduBXF51zbhQgiBAM/dn2PwqQJOxsEcNLlW2pTpPL7ehROoBuj8qwEP3B
mqD+MLheIEOvXqPr7QfnHhKAGlHDE8bdwSGb5OCj5hNY/WzMpyQiD2ojQGapQpVn
UodXA1oDca9f431rUv0UF5ZVgzKE+qmhaLuNNMAs7gsY7Q/+c2ZYWnpOX1yu8Zlc
1yXHu1FtRBDt7FicI8kQvBmVMQApepnnbW09HMbB1Rs5r+HNElCKUpKLwHzDzdyc
0siasC3XVVaFHVWqcGZcHzvIsHP4Ix6eQp4pRUV1BvLXGcFI398mMWnhSjAMUR4r
urlcoBEwlAhI72ScdYjj/T3rHPo2T2ycsbZMHtieKEO5OiyIPYURZxKiBtCHdHM0
H/4qACnaYdwf6ukea3RC/R2TxKNN9U8m4LSDnmFEBQNKSpUtOYrHS4K8HhvQj5mN
jTgwmCMSf8uj9ak16YzT9WSubb2tAygvgSzwpyVoiWBH+yacUZeP2x28V24WS/ZA
2Ddn56QCLec/3p/Me9006b6+/xBS970v+iLuCzKDZrgmIZ4btQbJ3c6XyN9hGXpc
rHAgZwK/RIHqeRV264I+tpHxYDxtKJIg57fV0GRGHbe/suMWOBSgtISsGfJ9XwGn
YZ/uqEBSs+nfnekiZSsJ7iclu/j8P60bF6WoSEedoAWP/J0tmB3rvI05oAX12TBA
4tk1sY2L1/6O2egqfvX5M2XFYXMxctSz/kXKqGvuoMC2qUYLqzafTnlZ4VgZNz5p
unzlWPDmfalUCGW9Sdz6CYcJz2vsBm8rvwkm65hJ5NPueHehQcxBPCfqeqVqwJ0k
bfTi7RefLJBfPu9+2JS/NvpgCaBgejzWnocwb90DxoLw6jKdFDX+ddy42el/Ajui
bkrddCqLxZguyg3CymNlXph5UEuf679h2XVFPHg5OiNTMZmwV+Jp4tnykvwbXnTG
aMybVJxhyemOk80ucdAphfarVx2JD9MDdaw+VJUWY+EGKnFTKX8b77zZGz8Up9mj
G4dF4JvWa5D8+HLNMNvH4cyjQRvb9d6ePKw7elVTULL3t68XIKZqicQb6A6DTaZo
tN5CAMqRjvdxV9uKtjlsEm4s7amQM8inxjtMq69a2gi0dvmqcvnVM/0oRDCbs38j
y1jGb2bpXkzR6eaXTkMoLe9Dp8TWmDXONhctTMusDPQIhXd2SWHWg2QF6mi+dO0Z
FIGg48MdlcrLXdQZsX4+/Wa7pALUbqMzoajygONlfWv9iOY7ENHB1ZXp/p5yaNMu
CoLCYxoxdMW2TB0LQfLAYbGmcWEROLJnxpZc4vfaePKsDKfSgw0N2xMFbalxQiUv
JxWazKDY70rz2AAGGX8qkQEHazKIJCJwwmdVCRIuUQejDjMCC9gv3Q4T6eETGkfh
xA+eaoS0pGn1hilMuYVzQJfNdoh4ss7Oy2QvVpYWv+Q826SPG2UfG3CGN+WhK/kB
c7JYA+ZTiFPOfkFJ0O9j3Kaqn+A0G9xfgQQHj2FQTXWXw64tv6ZlWmvcU2ztwOTQ
WhyrMTLkLrfiO9YjqGYzklOzrqQwlhRMpvKDOk8s/HVegpeQ+nDS0+tZ0oPaofVz
CP4BgxjH8kVe/DVYFYgKqEFgZiFRp67XH5UGjCJWri5lbQoEjrn1DO/O5H5vAubZ
ndk4HkFsdbh/xTNAhIs4+VExGjS1PlyPGFlJMFx0wHm3h8p5dTR7zsiJLQwdfTJp
rmz4hTEiBxrRIaygq9taVftoCRc6Hd0f89jtCyUYE94IF3PxbAz3twlanL7TqIef
fHOPcqljUDW+SRZQpcR9uzZhq/fuMv5T0dn183mkZh6Ya5c/zW19ERjUFnWKM/0m
NboWP/tIdtERSVEIGNRKSUsyYZkqD9+aGA5PQlniR1vqeKDhIfUChueW/iV6QZdf
d4E+XJqGMaI2TYUJN2yIFGHX4i0hP3hD6bBrrngg/oi2czzbvpIJhvlkzp41h3Ky
UyICp9UQtncep9iOTtpzpLtYcjJumJGmSEeAZdMoaog4+wikJ0TSuDXvMmENdPqx
Gtsw/xIjEklFoYGNDR7ZAaMbloIxMRxX5uJSMrmfqcnPzk2kpIJKaEVNnGy2N+sC
AOmfsRSrCxrDYvXELpii+FXyc7nyfUtudGLxbeF4aLqNFT04vVFJoPFNxOLXRh2J
QQYX4Tllf53MQMgpq38mcYn7uqUGB+Wppj9YedmK8V+fUbl01UUEnUGMAUkfPk3p
zmOBIJ0bbc2zshbPBqiZjrbj66Hl0YxtXMJDewe6ekRUTYwhghJzDyj7hSKITdmr
zFWln9rWG5JJI8yVlzM+JeO+GEqBy4Px++RbgqPLd/UxZ7R0Sau3GR9l/GVz2x3/
RDTmeJvntEs6XfC0ntDQaCrQbnMIUJwuiQGXyaCYJmj80mJ4zj/yxWZv2YEqT8F9
5gw0JkxActCMAcz0j4TOmydhUCIj5CxdKDM5O3PToqKNrWp4D6+UU07KWDt4nZsi
0GjecShQgshYoXGXVr+4bPta+xWvz+A0C/3n9m6DF+Mhnmy/QOLF1rjP/gOFalsg
hCXihfF+MbSixEi87T11mVyMF4UocFSiUO1+AyAvDydZwpwuccQb0CLLSY1e4ulR
86OKy6PFCRT8k+rUTRD5dCSqbdFtnhkSYCMSwZos0pBWJhaOWLwQnjgA/C8GIkP9
FEqhfj2ACgGw3ddTwkA7yr5iORkxIxafax5n9NUsnDXwN/Q82ZIlK4Uwf66Wj9zV
HW0oFjlIIWYqxrwnmVDXedH2cF+mIWh3MimmeER9Aag+yp5jmftaCDZf9pcp6+bj
njhBfxvevMK/GiLIJMSijZAyICrPhpzj8reduUjiBULnTLY0jckCpY8/vgAuozwb
lMDKInDn3kfAfMJ1F1ir1gShSItnKodpfyjJtf6vQpzuYwdB6fRFeOgIskJ+GD3s
R2tXzXAsOrkf4r5FlaBbt+IKGLyx+Ewdqz0S53ewt4qw8KiKN7RUKqU5nJH4+LQR
naR0zbpSyoHpalwA5dDJ95GDDO1t7H1dJ262utNzpIsBF1kb2p8jW9VhA/svUBI5
uutK6t/W1PKRh80Wnqa2zQfsNCRsRNQhWOyxdC6h0r92+7TQszfvPX3eEm3OpDfG
o7Bp8N0JJHOpiDKveNwrx+ZtVrw/TxWXahI1BNxajrdaeigIHrzcRahD4fEmFox+
pNRPM1pAGVY1f22bAmCV6asuA+T9WmnSkk4NJtQW+ob5c25Z8pjjovDRuC9rRb5t
9cUOP0kONO6Ylgvn0JsX9REKcm+evQExQWuE3rqolzsyDaND14Rcu3DEQCU/6v6Y
BTsBnAiDCqXSKIOTwq4tzAKK+iKCrBAjYZEeXLN9j0e/w0gCpkKKL/nbe4jcShjY
NmUwI5/WcyRm2Lrj+/Ymx8CPwTsove0yUjf/+WAyZ95YuwMEpgejSQUNJU1XDDcF
rVurMLiFufvap+9bhmBoOzGbMIcy+lvAg3Ho6lXZy/aj/jKN39I1WFSDJc4+rdYO
O1VdDFDXh3FRRkhbeJbfrwVjvjvJO5/4bHRxlJuiajgbc6oop1sTtVIC+lxXL7wn
9XR9BvaGihwpx0n1t2i3jtmqYMcpHuqfFQeSSCR35TdcgauI3EPswKQoQBi95qYc
9bqX+CfvjNdOBif4xglzaJlTeoXGT10YfNjnflipZoXa/RFzDswLA6m2CNhnhA0n
9bTJfDO1wffjQNUC3o0+AO4ttsUR2KT45k8u0G9NmX8P+4WNKQb4I1Cf4HD9ZTHj
FMXGyEeN7l6uKGdlH5pDkC6B3ONfACUTh0+cyemtVDENXiZYUwQQVdh1q5CQpVQm
dkHLxkJ1C9bP302MZYECrqLzFbKjtzpw4F1xuqy1zorrcuKvPiiDWUU+eYY0anAy
zelDcyaKwuN/BfAoeN9WNhTVQJ5rtKXtdhvbDXKjowPauCj/IZOCr4ROYgz5XBY6
0yz7PfEl23N9sPq5F2vQ02ZFZYIfHXthxLfm6HxU3cV2YpFCvNLjRahsuyeDtPKv
P5AhNWYXw5O/XLQeWS/t72zT1ND43nVQ7QkZl7CJ+2qkprYBwMZdbwkz9fsdofkQ
Nw/GWOFzb9nA+AZpT3lyO+VlO/s05ETkiNhCxapny54AobxSTM8BvmAUHcqyGEBH
ipOKXZCuEZZLFL5drrbi7F1aJzq+inKjvkR9ihVDxbJq0LimwMrmqvovCoEkeXUe
rAZ6Wdqxzvf+oShZLV6639A8Y8EB1M3Zql0oEUMk6iJBo9tlN3FjDYStw711XMUP
CzRguJwSRARxeL6gfsWW+fC5ekm2+SFDMQpYZuno8kwPgAyUFC1NABdGbkwf5c3m
O49/Gl4L8dfy6fbfJ1+XygrqMieC65g/+Nf+m5HDnVu1WBFu9QjHpWbjLGTiZCCJ
82AXi/q9tkewAOUJia/uMTmgUZw4RguxdpDGHw3ISSvCI1YKIqU8zoko+0VUtx6S
AmokSTa0UT45ODk5Fe/YDBfi4gI+S2IZINzILyLRFaAjIvNMi+P014REdccyadlY
xXwGh3Sl02olbwScjkFCEAXa0hLoE8ZAfh1cbgXdY4OgMuEtXdRiyIVOfZJ0Qs6r
Kc7VaSMnZC1fEiZysedBRPl6gmcl4JoEKnw0QjmAqJKVuSBFxbc0fmkUPUPpMXN5
ZXQxTxlXY8xXUnnggQpWLsctnIse3C5VlhvqZDVNrX/gBc8YH/U8ONSnjGVsq2Uh
sRJSSeWrsYHYZCC6EREqjgk3JRlM7co19D4WZhIelO6kNRVdIIClpVvGFCMujX2w
eC3BKFSBFqE1FvEgO3uY11eyfvPUC37o5aTHnmBaWTDaRc8KbYCC6Tqs0phSfky0
sFgnWNtsl0vNLZEOKFbimTFCakSn8xUTd22pwe8v6pfn3PptTpzslpQ/70qubyN8
fsX9xv3CqWRvzzfepCZQr35kNc0mCHp9I8B8n3k5+TV4IgDfWK/6m88F6pV418bd
SqH0yx4hvl5xvHStDSxgFmUKAD46DWnJuK7GFXseqNrTu5yUznajLFDgv5XURfoD
SJP2mng68raXaZZhxRObSCDxpTkH7IXAR6Yrp6LtDuIHtxwyBfRE7EgvO3YQKn6M
jg3YHMa5yZg+6aBNycMIkrVav404YkzUtWbFait9h/HudcpGnM0I3w9ZERLlLHFN
FCV/QYP7Y5/NtKxIizzsCXEHnZBGGH80h0ilCt333C0+a/RTkooY0NKp4sGPOdVI
PHJ7qks/wRzeRmqpBvQ6eohGTmq6D95q7J/QwXaD/iaDh+h9MOZW2oNQVS0TdSbi
BgIyIpp/XZVWamFI41moSSyUmnfzRHB47nN/7DgLBV8VUYT5ICeHnehCVvSAL+PL
i4Tmfjzg6AxISvq9f2wl5zkxFtUQyA2ASlqhyC30DKHGLl2q27TQRMajbeTQudes
zzeCMSaMP2Pj0quYNYS8DPUhv6/QO51eLupg1eRX8GF9cKu8Z/oqqn9Ly/zeWhzz
1wFgT56LjvJafjQWwXvfdLSBrYJPAYpw0NZmF+FHWLkfr3eA2gGNKo2cEHjhRg8U
ypcBq3xb9OmkDP/G9LTHjORlI4Bi5jGFj0hixl0mHvdhU0PW4oO1AJ5J04kc0Ocz
k6pwiDqZosA7j+pmPOfC9TRRDsWEWbWks5xPqqdTekLX3WMqr31Cu447c5q8/jD+
2MskBn261VZOAhJi174OLSao0hYKPmx2vxpbpZzgznGOIWlogyoVYP/LeuBHcRH7
/NBoN7rJnSD0DSrV0E0+zJJcswstFbdn8X7x3KWekfx8KgAVQSMbjTDJ6nR5Jz96
PetCBBDstgt7ki7qLDbtSRgWSLzj/dK6qIXECKXMFf1t9qH8iLYK4gcXuJC7Ihak
iUkYPk/bt3jf4V7nJ9QLu1Ww48GGjI+DYE9DGP30oJ7anxjxr3WcRZ6jUgu8TODQ
HBy8FuXAIXXF1jNQYYB/lCNIGFPEyPtdkoLspRVbH1yB8YYAdKuZoVJqpBol3n/S
IXMmtyW9Fu07ItndLHdA2TrFfiXyQ76i36+IUnjeSHcRo+7KJm3V2H6uAxVPvnbo
FZ1BtAgdYcGFxaaS/azEat3Gnydd1Mk1gRfh5d7qYVJoJ74CilS7KqscoTEd3Ccv
7Wj0L8o4GTzqlxmzqu42lY2r9yMWT+OyBhs0PFhGBAoQihqcuA52pyb7cqPImlE8
FSBoaNhhj+2jP/oi2+jOlZX+UgID0XW5+pEAgg9TZ3D/MkeZlCKPC1mWeeGDRjFS
Vp+2dXiTihuVDGEMOoSdBwOFtlyt30T3fpesuz/sYzEO+XYCmHZ1+90gfmm0ZYsB
+0j+UI21Kz9gXU/Vb6Gl4DHc2NpZMkWltaUkrau0IHdjUWvMU7f64ZjQxulUek4M
NsrQX2JpOTX7sW9r3zf6EWmWCRjDVXeIysqCQIgSNSVfoU236xJ2/n0PmPEdttip
+ouEVvE+jvRlMtmv9x25FXlTYnO/LdLpxY6vttUa5PLR93dEEgs+Pvv5HnAcRq+O
/QIzpxt1fAIA/Zm56qG2AhUWtWHNhdKeG4mM1c2xyNa8KXr7fAQLQh6bjpwYYDYL
ChQd9zgfTvmKbN7W4Amb+FBKVBbCsCk/zdLz5dGbGilSqaLzP2CcSLxxXHwjaeKK
ZMxFk8MJ0gW+xKFef+z1UxKHzDBxNIM+sw6fl/x0wQr7GuQFjQxB7Uutw4hpk9xy
uW9S1uXYU9dyXQfqkl3Iax2wFLEi4My2JOgHxsvftEeeF7D2yLzrxpDuXBBEdsjU
LQCT18Je15t4nAs46x4n5WNlZEd0xzO+Vto9KEWykRKRCMy9xwb8tHE5KmEWu3yu
T2zOjeCRoMpG5Y/hTwwpT4uz6xJO05aYJus4WmXHLr8TGQfJ3QRh/9zweqOYkheq
w/6vsnjgQasejDlAyjbvIAjZqOEAXvGMIDoRQ+U7ydG0UCq6dhBB4HvQM+pi1eCt
+5186DpHWbRcnA93Ig44p2xtFBdN+Y1MJXTW75KM4UsUU1gs9T7tOsvvG3AJ5X4L
7BZultDcjJ/kB253vUWR1wqvgTprdhqNNo/NdN2J2+0nheSs86PVIzUaF1xMELsr
iBFTUYfor9OBKyVXihgmIxBxnoKtgB/75AdZhttyqGZFLqM0MCUayFk3SKon8lrc
vLxlq9vsYXeTASeLIXAbRmrbcRNePF4tn1bmDyZ8+2GCOFr7j0Mwp6SS08MbQ8BJ
tc5IEKa4YJ9lVLjsr9tjnnVhpGijvp6nL8tUoaPZkeQuVv7pFWUH5LKNEWHmsl/Q
DVlOwGVltQ7k5qPT1vUvmXeCbN3xp+wI3LBpXUs3tWnuRRmfBKXKcFnept8b4OJj
/nMwqwXKmWb4JeMN3KbjraVQgz2rrYCxsCxmcG184ooUEEA5khLdlzf6cXy4JSGH
EeRzx7FUaTcfHuOi7VjoMu1TBBf3ZaAzbyzlC2otL8DoNAwA+ptkL001RmQTo5+U
fALn344X/9sEngPUURhC6kqaWfIyEGZDDTPOObXbPjLLvalTKIH+SsnNEN73RpNW
dzj8jNexJyPc7AgzuCC9Blz0VIQyUXqEP7yFhfBB5ZG253y7dQayBEQIRNX1ahbc
917/Lr7Yf4I9II3YKNY4+gpnHw7VFO81cQfE3jC8re9ZCYUa2qJWY3kjOPSqjPfj
W1ZatkSKo15MZUrIn4ocLGxppQ1bXGP2JLFp5uwVMIEbkeJUV5RPPj8FL/PPnEMr
ek2gm2dUnqIth5S+q60rNZncieDXbOq9dCCYwIMp/sQBSYJSwUw0kqJaMdUCqr/U
YYs7+GR7HpmeZVhpxflqEuCispT+lMHnNLJuwLS2swXt6hHyx6kO7edcPqU96OSp
xBRtNaCATnm2xlewnJMa6ZVIgyBUp9VHRAA/aqqWU5HrGUgr/rLAj8/zy+CrHj79
QvMajiRkcO0qx3vGkPe6G29gA9UyTwlq4Puh0mdKSlj7G8JGVaHn8p9PF1RIyPN1
NRWuVEjtiEkVGKwYEYgAIn+wkZS1jZy49pg1IiU8FIXbgHQm1YT1IGR+4V3slxaz
45Jwx6Ei80dO0OIXKB7GK1TMp0dp5S/B6HnvVUaOXIx2t7FOAuWtT7Zz0SjvbAtt
usVLf0TEk7OjbIc+bKYUnENrY44aYOw3mWlTIddZ68xs2Sh4NxZHES590fdbnnBx
QSMsKP15I4dnzW4YPL1+j0gfscA9Vaijr42CeqJtbAmUjcZe8nsaSiIufLE4q9kJ
FmLXm/TJU0hdSs8y/0tICzwSvraX4vFlln7UJ9e6W4jXEBtlQhwC/9Lnp9h3oUKk
q+t63G3gqhvq4YB5MVnpmYQ6mmUvWWW4EscjSA/RIg3SUcP/5uMbDNYsn+JYF6CS
PfJfqk9yWnVFve4BbRF8gn+y5cZwRT9sXFdHV8NHkbRotBB37AmTUBFvMVYziSSu
yTb/GQc7iQXTjCN0PbopYakydcVs6LDNny1s6gNYC3ku8NAnHhaef3k033tYYEXH
UA2+4ieUINUSLAhmm5vgH+hBaCQtzajhOa7AYySr54JwxbqelsRxqDW1rUgPxq55
IMP0Wvt3EfUtBPVyUXi4wyRuzvmYbgRfx3kz/N+51p9q4HRVhnlML2wH5pLTRL5G
igoRfInuNLgIzW1SGi4eygEYjOLNuKNg6pIbumwj1kOKh+RtGgWe8sHnWxNRorfg
4SN3a1lwBYG8crKqCnYpcYEMzTRPRJNcvV5AF8ZaJum7gfJM/fIacnXjj6TllvoH
Et44MiK7LP+n0zE6GAEL9LNuEyjyDhPZ8a6Lvr56ybbgTe1FE7eZEjdiWIKPBzJH
RB/PIZ80gwhW21mhf/8gffN9z1OXM1UhPa4lRb7bx+VrRYh1wmjydITseQuOI05a
FxB8t8ARYkgGj1XAeH4oFA0YnDnOsyrgdiahWd1iloIo15jllBIKaLbc7FCrEKsF
Trmd94H7JlAWeiHFhIQzT/eOax3vYc7ORjU0YmUzUh+yqOIKohHbEqLi2K0lZFu1
yhinO/yhmWs1EFwH95RVvu1ZrPAmUTJv52wAocBXHXB8bo4bXjJmcwyZMYs0qB5T
ziJJdLaZuHHUFqVCJW740tZWr/YgK+zifdrfHlNhr9UWWlUVUr1BhSFx3H5Vfn/N
far3BASMJgf2mGIulCENLdQTr7JdNgiS4VHcMB0NGkNb5jAGd0GP09PidC989tbq
3aQvhQY4NrwRfjZT8PtoxnZZUt36Sgf8B1pshzTEYAwxTt10rULOLWAD4F5hIVXv
cWeLcUXGOahHGVKKevnicus9cY/fGFMjj+ubekFhy3PQjS6rbBqv0q3RVcgS5Wv4
i6gsNjR3yfa+twImKTmRVJQSvFhJZ32eDSYl9CGnrntavKBJR/t/mr4G+lJZ0CUV
lkr2+0yF1osLa4kuvWBvD/ujHNssziAzdsarolBQeluNKIOMBuN4/J0RNPcl7LVn
vXVu0JzUpBXQ3AooD6DBDFvffvqHMYYzchT8zgHsaIU+HjjDB7xQtYj5+DLSz16Z
4z3HF0whjNyV14sC2ebWOgL+51LO7Amo7JlEgcq8tvWrTLSue3l9ZTcclfWkRWI9
nBTBTSLQFl+NElMcuJXgou9LWpEmuKX1AbtpIokXlDp3/zI7KCZhxX0TRGXGm9fe
w7FGm5Qd5WDb204hj7dynw/9/hyv9t783ECcjS45z3L9jbo77S5JMyR+vqcz1jng
eTG0zdslXWitCQIfyFtqFXDpYdAF80v3k9QWNV3B3zuinYV6InM4s0x0CBNDvZ+h
BLUcvIu3h071m8q1ts5Kr+cLR17Pa7rwaP7kYrAnKWuQvq5ZG7VzmzQRz+avahO8
tuOxlgITXHBUnmDA+n26VHOW4GflEH7RPJyU+g+nTajaYX+9e/rBwQGbHF/rtGS7
XfKNpXsyUQp+jbTBr8HLlZKGS6s29IOYDpqR/Ef0h6YPakix+txgOiGTKevF9Ha7
t+8C+YFY0OMYi7wb0NGMegHn3nJ3QB74JnFvgHDBWmdTniocvW5w4OsX1fGoonD2
2HYIxHQX0OMf9VxlD4QanAkQ8B9D3hCon5fUqC3XFet1Mi5EdI91XM3MBX6A/JlH
uZUC87yZ9TkYKm9YE1Ks1JkLIpnd5xtY3Rurzy7RuTPDjwTzCj6AXPIEEpJRfBCK
EZIB4vqgvRCxWwsZkIVA6+Lzr1TSMhBUuLVjGq2uGmonUwYBgLp7ogOZd6VzXF+4
SGQPSff74y4cHNdz5dK7b7Gp4aDvMjeYPfa5806FkDgxtdgsGzAcfnx6rPsUi6yg
Xi/15j+Gaykn1e92GhJeypJ5A2CQH2ENS6Px8NX9iAQiFps1eTBpQ8C43ifxpcb0
8hgRdddPTwHN3FcdnYNy3LtiIZ/CHxmgRtuuQ8nGdajSojIWi1WUac9YfHe7Exn/
x1Vbson4FmsZZo42cK6rZcwRg1tEr0ajqQh6J4oJi0ixRP194u82ybYXe0MaEyia
xSajKXKL1dTEn6pBnND3D1R+dz7ZHtZsWtCrGAebcQmwVOc2qt0ybtX6sd0Lp2XK
uqVUBfJp4JiGpjNMLW3yPjEiKT9Eriy/k8zLwqoXLe2BxOVcheBYWiVGNmoHCWqL
jRaWfd6bYlOoYEjGj9SUMHGqSLLxYjEgBE0hnyt44nBhfVDCEOaV66b3tltR/4lt
Nj/a2wacjZtDyJvQd6kBr2xcKSvBrc9qUJUlObx0Z2QBdLY/BRb6nFPH0OdwtEyF
P8X79aTiGrGHoZBmC8d8+31idd+k/om+lx+RATm1UruS0d083vKly9Vg6c8OPpOv
f+zl/gM4zpuiyGe9hxQuZUfv/nSiGecrxFfOp3RLcHB3G3GRL4pYc9SvKM1dpsUb
7aHJ8zqK+uDE976C9Up9wUcqpbkdkcUrYdnFm/PZ+tsWVoTRd8wejgvk2tdarlF0
HZ1afCLSuLua7xtaRtzkfYel72d5+U7A2szf+7SvLV2rzfFI7ghKZWk5Jwz/GUpE
9qYqgpSE7YaDmxDrfYw6AqptqDdOI4ocdAkTiQ1TN9WTcPjQQZMFvW75MBzCXDgq
zD7Jls+hKvpjMV/BLPgYtxGUFjNr8z7o40zzOVsvDPM88EP0DOSLjvFeS3weH7us
LKvnUcizxmpcgICNPFqgvlDMn5dLbP+Wc4O/ABdH+ZsskAuMI/dYC1dTP09YOmBu
6pYS4YAY1u1f0IXOo0wbr7djcW7tlbWBi4s/lck0mqYtzoaSUSLvqM0elf/DMzv2
3VUNTDTe932wlMSBLfXSqC7hI5B3htGLKPLjKHxvxlgo2rPppUYrKaaU6WAWZs/O
J5UNdmDnDBJTwyyDQI5cYrsV0teZJlrPOj2zkRlM2iXIKgEUCDP7eG/H8dWycfxq
9FCQKCuvSgvpJlK5/cFC6woQBNu0F4PJSzAht3XpWlSfosPEOTTqJZi4buMVx4/U
MYRVL2lMpv6GTYG5C7YzOf89yZFdX4bvLScYsEjDqLSlZr5Wm4xsQhBWr5q9QsP5
C5uDn1RKdFyThMT9GVh+9vHtLs3n2fiPgBtLaVEBsIaiioqA1jPlVLVcud3R73TA
UxBnFYhDP6LvFXouzocqeVgDMMte+3Lnkas+CcjONgq8AW0aZY9IamSV52vHWKBc
fAgTeDP+n7yraqJb0/uOzfgvndXZPu4NpSs+jHE7PsgxKt7uZtVQwUq9guYpWZvh
wZg/d6rP3tw0BDkPEI4g6b2VrBH0H6VjsF+FpWo+6rFv26jT1WltIxF09hbG4aNc
B6kgidPA0WTMS/D37ezasz0LAu5o5VnjZ84jBlkUcW/PAFBFxFlpDfFSK5ynn5SX
bdtWAxkvqIe6OfcKqEnBy1mKf/6g9+7PgfGOhiT8JlWej3tePYnVkJaNPW6QGI0k
5ETzfLY16nAzE4ffXHPobVejLsJVjd+8J1PtjVXOabSW8hY3U2migUwCMf6uX4qK
dp1dsVm067FqYd+rimkoOJVifIn9Du/XPJYGpGJo9zE2unPKiu8CZI9ERU7JP2ca
l19NrdCo73D+fhXdEs7MeiNjkeMfxkp3WkEGAO2uF1L0RnDaiRrD28s4zdjbT6C4
B8weYYvx2bQ8ndNIdYCjn2fsjGj+Y+pgGvS/zP22zikol6ehwqQNv39RKQ29PH4D
U5DTcTjax3Gm7Lil+pmDRmKUq7ePi08caQFsDG6e6BBWla40jtf0kV9TGNxTstyo
OooVW4XcL+WzBu6YytaSv8onn0i8mgMFlXc58bSQIewYwkbgRGjwQe5J6Y3kcMtD
k/hOuDHIRBmknyo/5ysYNxge3x6s3zSTlVQlNbwl9lmRzPR1+pAQC8RLY66Pgepm
2sui4nnO1H+qADrKMyMudXzm27mZN2QsvfBB7/Be2doHcmKJ3A+ira3sksXK3YGK
Y6QSTFzWG/c15nhjg6f2MGLwb4txCAh3x/R9feWj6aMAgdwvp7u6Bq66QAq1IKG8
lRsNFMRUAh9IPRDX8KFrRsPY/SfPrZK/aSbiO69tJkki14f7RHypTw02lcmr4d40
olfqP3Jrqp1Glv2cx490X4vsL1fFlJ5iwRRttbMHcPguJmsuWdvmzuTwkmhPshw7
15IxXXRlHQxyPYxdcmT14H9PO+dTaeloJrk1a47Gm3WZETd1ykjvNu6f06fMf/0Q
djlEIpGahtHeKuAAOqW7fl0AvY824qtof6h3AjRfmvbuVow2ci+Yea/odi3ac+R5
saTLl5TBr7gbLBIWv+zgWeeNyjrtSnGAOOw+BNRrWUJGNFuBuuyKP89U1NWPV2/a
pV5McYpVPtXH+saa7OWaq6toZFNXbsDARtT+KInrZ5io8jGy4om88bV9BMa4NCQ8
J8G09RUQVg4kwISnwxqWYMpU3K0sH+2eUgEFupxASv7f2kPhs0eB4FXb9SvLeuGM
4e5P83/7ddCDZ+GVHcIS9hhzUb281/qr1zLus3ZxHKReAZ94Ql/k2bWn5bthYFJQ
N28x7oZj0lU6nv7//XaYRr6QZih0tf+kVGAKOeOKacZyaW0JAaDMyRFjSb6IZrFr
PKf4VyDjDxLB9JCQxlpBHk5akR3boZ8dMstWjB/wog6mLQb8fXAdBF60xdRu+NHA
zNaNQJgt9P6TL8Gqreeugz9kZlP/aOCeTTTsWweSM+hyWXZzBUgFSE73BQUDzETz
fROv7RyvbrO+jusxvrI42UmIEVtGOaqgOoWYoC5l7vkEx96e82UnKdHcOQ9QIVWe
egXEYXdyv/NnR2DNVCGE96v+qVBPXcvXPCQmd4yX+5ApNx8o/tgOj4YLMh4OZUP3
EUDhRhVv47ehRfzxaHnn/qO8NHqiNE4acACJ/BVlOF2GgQ7tShPZqh3TEIZHyapM
kg1V0YFm0C9BEULRAPrH2RCg3L3r+xNKkg0r2+GpGmIRejypuofCqVCAzvlVvlq+
8ist2XY2o9SuSnLiHH6cB36a7eoLsRSitWFalQUkwssvdaPrbISksua8FbvCzV0j
eDTdtOENrDgHuhOiQQoqA6tMLTNG1F24XtNHlmlCCasw9dMw6zdSuB962Z5sZFs9
/UaPWpVoJEpXrr86UUaNQZzXZ+j81Cs1d3nnculecvDn4C7ePVC+i8FfieZNqnIa
GNNQHrvEx4uRJCwkJEyy8xOOZrWYjAUPooY3O049zj+PxXLACPhtYIKTDJQOTNB8
wVFauuQPPf+C8An2M0uptL4s1CtpasNeCAi7HpmWmS4dBIgGJSL2S1VC6DIuoCwG
k/FUmKqjA/kTJGWzzaEbAzGor7HVchkOmrOmHQ9fKSWGoOgY9mzHi6WfEZLwd7zF
opN66IUcLa6GBxlpNh8ibzFWhzuBhrjzyT4UDbYXTNayQKsLLle3Poo2HK6qnUwE
PmTB6oeSI7Ep4kuMRy8FawLMCVin39rKOMUgS9t+1tRcFHUB3Ak5heRlvfB/5WZE
Hg21/RTCGP07nmIfp75Uh1ZJx44JThAwm5lgPda5dyQ4p67JdWxe+5OyS/Vcl4eF
7aBOe727RA++WM6V3JVrBGkQKqFvN5CU8U5Ymb7tSyQFYSZpVU1iEZqPi72n4Zg4
JcZuhcnDetKHGH/NgkpWD950o6jmifqQhsqKOSkbhTSyJMxPHET/54o/CrfbWgb8
UdZv5QK6LOB5zOyKzkMz3ovuRdCDpEhDefqK7JhTkdleNNUJKkNV5tsH93b0K0Wz
/ycAFAMI3Tbt3DwDq/U0lUhYSrHqA+LkrZ/n+czZU5qFs3ZeTjDm2/CoaMFYCem/
T/knsszuMJQlJlc49QoZB7YNn2lhNQm3/nbilH+jQzG6oRKIWiySxGE/Lm4fFgLa
Ul+vQtDvoonhiliwTS2psJPX7uJu7/P1R8cUSfb+OPghe4qIyhf2FpWEFSCn1iL0
cAakrL+0zde6pxhsNunQ+ueXQ2Xl/9IHuCn+uCpBGzjL2trcMwQXyvBpjx72N3jw
TUKPyRUXh2IHrjEOGq9vGoyIUJHPH3uUHFzgmENKLR/GXu1lhFNkJhDxzbfls/V4
6opbHrJR9I27eDl0gJZ+ThQI2TyNa2rPn8zU02NaA5LlCXMNQuiBmiXjFcXL96xB
DnOdKkC0URO9a9zOmznBma9QodPyI7a1Z4F9zg4qowfyLXoqdLpkTWG5hfQDNf4w
1jdf7BFNKMItGshB9puVKKQJ6LuAbG+kPB3jOxGloRIG96LDR8R2QvY8i6xo60dv
Gl40GrJpgSVdj+oawnCDm06Sv3zKzU6SBtO4DFUnMKrRV106at3LVDfvmjRCnd+5
OEGmztbYtYC4MWy47awYy9+I7yJ3TP+kWgR82c8pWg3QSA1plUaXJvV6hsq34JSE
ol79p3Y7Z8en68prutGwqZ76fWXZ9VFVc6Z2kxLnOBzLfasqKqnUy5rBBAopocrG
SOrojbdgooKBuRpzLCW4dnjQKbESYEW9K3FJNUtSKnp3oFu/2uH4dn0VnGQzIHGN
DAp6XVZ5OT6GH/cjpFfixy2hMGdxDQUz91O1uiyYJfb4D52y3/hOGYUfPlnXRlsI
c1MjHbH9Vqgd6l+XQJeg5GMsTFnoMZ/9hCainlTHTNsRt9lg4XFCD9DzUA6ebW5i
F+uOTF2SAsYNcjAqHl2JUTM3thVnQaL07X5S2UXH6uB7fIbQOZtFgT/Os5x40s71
A7BV1axEh/jYyFQAb7BRXWBVdcH2P2eMjt6HmRYu49DDdBRWLj+9AyAC3PCOiZmk
Ummn5bPFP0QT/lB+L9Xc0OaS2faYm1+O+ZExGSLL9twUQDuA0YOSOTjc6L32a/KV
mElLZEjNkHObIkZK+sxebTNUbEkMc+dyBnKjVaOsv3JTyF35evEou0Ucd+OtOVl2
TFrMwyq+Y5s9bvmz/6EMEyWh5OmjhwDePPT3M3Bnq2P103BrWYxnj9rql2BHJ1Lh
Y6PrYb9l4IdezTXx14vp9wMICOs9K9QjfpqgZLX1ImWmo+09MYX59tuV9Vd7xXql
2X85BRTPYpul1khISUx1UP/QRzZWtYudf3JdWoYmHp82i1HNlAf8qidqT/qOquac
iUlFy4yyTDJnfd40g2/ykWdmcVzLkgGt7GOaSrotT2lzFUUzIclsj8YgrzNlJXNl
ImujuCg5s4uuBPmqfiKK6PVUe943FIzf0E3feqrM6rHIuaX0U90LAquckmjDReD5
81vqjouD5ef152fa4zkx6bgJFEQr8001zk4sce0MojY5R9cuZ618LgWSI/S1sVnI
lwrgKE3bIEtyCFrxI+yywBXPD5fQqfZsiSwnrWbixo+P/UbORhRjUjLXQG0pZltt
9npjDVAsV0iBHTEOt/mPstIv1i8Z6nXjXEg0SrKVSP2hGtrok9AHhLSStcvbBqo+
pT1c/E3shKifZH1rQlrCDvu2o7s4YormDjeZbZ3xxwWuQbqSWsa/1DaWi3HjZ0yV
vXglENHLm2aAyf42o2iKB3UiiyE8Ff2rL7y4nos79s22bJJzQzzxfN4jXBFKm6GP
Ntu3W+MVoyJ3/cCHHakpKMBrqBpW3r8EXQI9jRgJ3P4mvKALWdx2vzDDOM8EtI3Q
+gENEgZ5yqdm1Cmj9AEMODRWvn0hkVFSHUFNlzoc0LKBS6KJ2ow0clFGIbrQXiCZ
v+xRO3ye1Qmimhllq6tqIN/LewBPd36w4PUsqeq9ywZiDHrbP/l8RLbM9kzIX38O
ih7VW8//ck3gun6h2LaLdmbBi+Y0v6iIorPXJg4JQK1Sy7gN6bl5BzZb97phTBXU
BupGOPaL8lCqo1rPz8U4Ne5BUtCJuyY63vEnTX6A/i0M7sew8V6mmdJHHgTGF4B4
4pZ5W4eh4AIY8Unhe75FzhP/54Kru6zoS8d5wxcyD2WtbB+2rAMBcSlIY1rHV2cB
OlK231DEcl0WOIEn9Jwg4F/4WgFCdO2Uggk1IMbqsUmmA1nLWCXA7Xyx42EPltwO
lMBsyz6mx32QzvhJtUeWarKQed4v5IfYcU1bCvSfJImNqQ4hJwXSGbOQJOsIWp2A
kf6Ff7gEUU10q3gyEBfT7/0L+hrqTcvNl5CF5bDJ7w20nZPkXPe8RJoonnspM8ka
nXWN3jZv36cw2Gn80G4VzcT8HxMHzi87XzTZXpSTRyWebvTOdFMc3tnst+hH5I6b
o5ub53cDV8v1cy5rnDdKK2iOj3mRq8BBfATY4Qs33DGGIlpDBaEcNPxrVMNfQsUz
PXl00GmtX1Ub0TDizKEHKegFYk4hNrV0h2NwsmVbhsCrSDm8nyYKQX+5HvwlQneI
Z9JxOYlPxW4kyipKxYVr+Q/D5OdGc9DAFRE+2gxiuXgGnDEwFygPL4j6Rp6S1PfV
bFLOSrmZs0BjMtAyq/dwXDxE1lDP6kgv4/8gnFnRBLr2DzFrel7u12jKIsgwsJQj
3IJndPqtYdt2I64mtq0U5mHCIz4RgWTZp1iO3u1P0qLKkBCw6sPu5Z8je4OmzBMs
AfMIuN5HA1CttWmqy1qQI/wdfmt1Pl/VJETrZXA/q83g471djGyxzJ8y4z/crLA+
q8FwbQpc7rpUtpbn9WHw3YdIV5V3VHFTG6Nw0tqgGTsLVCKMqRMyBRLBx5Apni+u
Dr07x+yz9tZK4KN8isl7APzeCbcx35b7gjLRWnX2hJkra/uSrHvCAiQeK9Q+FXRT
o3+WsgaP3RSHeFhP7EaazQSJgIU0Jn77UHQARbCV+xSDDSfXLED49gZo9mQHfdfi
fNB61LIPSFHzfbpLqW7C9qIRyewKoK5JWVfEfbf13mxhAW1s91pVvO9gUjhD33GS
DPSf/4wJi/+PicqGbBvAGuaYhcgGkG1KiXUZR8N54fPrrJHNCU4h+bGMpwbgiIMt
L+79KF7wmWineXO1VxVB20J3/1aZDpBw8RzNHA988jNVnrKljj6b1IgMX7lrGh7a
QygdUwEg6p+UwsYMHb5lCjuxC33vqW9vgaT5EA2ZXNausUMKwsS0/4WGM1pLz03h
BkqOfYVnB+PPCjojPiOmzUQfmc6GyjjZsT02pmL4gNUL+bMw06PDv2TLvnj5OtGj
gqu45m42VzqMHbHCXC5yCOODgY5VceAIJowFm5NqY4MNvZGibqfO/Op+3hzL5Z5T
jivmkT4ykeJemTBlbeF/FmtoYl+L+sqIHsIXtzkR11/Kc1WuO2VUNIGc75eWQV84
upAjzGiFeLJh5yJMBZ/B50R/rn1KpN1HZYUf4I+1qbBV60kCPfbkyuiMwuvX87zI
xYY19v75TP/yj+qq4C9wI8cmy/GJ9chkgQVhYgt65H6UQI9tR5dCrDysN4FQMrRu
xW791auxKqW6HgnpvrLa0SwdCzdzbIn+xRy0aR1NlATuPn9lrlvPc06h/gB+7+DG
PHeS7KqYYk7qZwJ/Z9Sf7CZ2vAzZvt+9UQxUVAHOafXe/jHzUQSA4JPhU9mq7Qca
qpXGZsv24uC1+SPVOZ9a2leBiGK2eB5ThF44QibyUdx4jnFKShsIA1zl2Jw7b1+h
fTNmT9tRlSvtvgcDgzIa7IYHdvXv4iy1BvqAwIIhYwSZx3TCSOoEz7atpBrv0K0S
FmB7NHGGGzV2eOhO/KK2l8S+I/3zSXqUWpvsl1fCnqQQW/dakDQwlyydyXD0DN8s
8953ZvSECzfEWY5QA+2s4ApZ8MMZ+PUQCbVJiUoqbhbxYMN39WmALey52iQpQYLL
Zb7ZqQevkmOlhl0K3sQTDRiV/JfQYN5y5XH/ggFWl9texUXzMcUAl868BH7vaRRG
5fGBy1V/0VL6eJhiaE93LSoSDaXZEmN68pvOw9+TI4ps4KmU+IomhTCGlhV/K6Jp
HvIaTeRTQep3uUD9yneYCBSB2HozAHalr62rIi+GWm5i4tUruKnZkase7D977vlX
zLEESWN/3RH14OnHxrMM+Rw/gJor9jlufNpSuUKiHsqHYtuVa72O8yYzmsfWAlpc
z3DSUa+3++8wv2Ap7IJ6f3I4nlzQZV/6MtDrARxv1p49PrmdU+DVhWKegx8gm9xn
kDz2FRLcrLB/r92OH4ucofA5Db3m0RMd7OEKZW4gg6XV7tcoFL1t2m0h/7TYkPqk
DrRkI0AIpg6V0qMCJME4xwAkNkymsNh5VP8ZW2sBHxg+of+oZeYxq2EZjZn2rDQo
zg10Zo53I5QL89E0kBzR0f7YRtA4Ig6zC/Vt765eVLkEWhYa/7GcW3d9VwjfSkCa
QvB8l4fmp+dpjD73ZPZeAXXXPdBX0dLJxz7D9CKYkfQJSd8fSUo913CXaBHxNFER
Q6dh5GRiHuxa4Gd1d7Pa4RsGnhRcRVJJJ1ecc3iX0FKh5bemyusb/ZZrSBGuLeCc
aNmsP6oH3YxL+htWppketOY4cDHJQU/uklA33rFQ+4TIUWZ4g/x3lCqPMFOcJG4K
0BM7KHU2zGKPtTr14d6hivwPuvyWBvaJK0q+GubbC4zUdXSAoOeoISEJbDHL1LJx
JJgsdnZccDKX+0ufusfIVYybMSc7bX9fRrFXPN+moQzaL9SgqOsLlkuw9jZY83Pw
8r73ibKgZkjYS1A9xp+i/0L+HvzlToefAiagd+x6cANG6H2mAsawlkBBC7mjmSwh
/pYqP+x2imU7aFauxTUeXPB04RkyD85Mhsu/vgc3WNJGd3/t7x8k1VTVtXqZf3ik
bx+LMmz7H8nqCpw52cFJ05CkiRMDhQ5mACKRvPM5Syyyt+FMWUHr6a/5vq0q+rft
ZYv4HDOkebOqSFrEHBbgdfq4QM1JFyjNufbEHW6T7VWWrVLYPpMt2qYPPdD6AT29
QUAxJzq+ddhKH3NnTP0Z0/IT6oaheTarkjNuF56TjkHsFD9frfzFsZOI7wNcWKMn
68Fyryox1sgSBwZUbczw6Iz4+72I3qm0F+gpcpUR5TYbGtWeu/PZONbksYN81+/e
PTXYjNiv9F2igqSD8XN9ZoXlVJnrsabhByi61NXvG3h/PgEcW9FdZ4apAuVCYMAG
boy10oJ+eVpKZrjOnBBhohsoYZTcZiwEMcShz+wDisfNo9tP8ebgVnj5QTRn1NPy
yCJeN0YDm0veEmctV0FWvkM/xmma6qKV5TCgULW3Gzp1Aei4k9wm+H/GdbBO9UDV
l9VSXNDKFICdzQIpwttSAy9ibb5aYRjUbsiI6oOHNRK6ljgcpDDuyNi3HcV1vtyF
mllIAiR2u8Kd5bIsg0s6lQ+ag4SX8Wsc+6tYWJEBqkVuhAGyZ0VJKxYKoLYoQeDz
zFUKvy9MG+o54tRyRKB3h8APDGWoUyMScXt4U547YrS+bzb6oibNtGFaElvjObEF
h2i6yShmy9vJQwf8X5zx5th9wyyggBqml5uwzsQKglT9V/XFG1gF/+5eqlLX4Qlm
ONKtbqt6y+CTtTqdegVMmkWEbHQUSs83KJAYB8t3GzmgHo0nx2FA1goIv0vaqjpf
EQEcMblea5/UJmp2eZD248WXCLwKGdaznhBr8fQ8XgiKNB3hnXa2HjUpxasQwUM0
vWNsA9HjbSkQbHCt6q+VH6bHMQZNrXwNhfFkFVfZvQXUJzXbMSxoZe8yW6W3o4gE
2g6UbgitD48pnBJq8pZm/fM2T0t/LTWUX0NxOxP2nO5fxW9j/FEnI2Kcp/oIStSe
Tr4LOi4/sXqZKGdrvrNjbwOhxiZSVSCetnUN3ULXcVoRLmj97HPmv2LhhCTNqCXv
BG3bumn7nAyFqM+FiFbut+K7tdZ3/VoLVBy96v7NR39Se9qvuKLsomlvm8heaeFA
ZZgdj7zp3tZNgkC/aWc2C49otWjAjl9aS32HFXYvGgPuk/+zhkD1mu9ntLbsbP+p
t+cnQVz5VjSnfeLf9scmhquj+tiEM8pmHPvPTNb6kEtnrEWTxrC0Gf/lgKtJArjV
+NKFaOuibu7m+wVT17TkJnOuEJyzN23tX6wZb8xqXAABAlRmpNVfZiwHHko7NMHY
g3O8BG2pDmc6Vow6hLcKt6OG+uR0E4yIvmLlsBhFCTWSk3TuVPHNr88P/D92pMoG
AUYRRsZv1toUEHpkY4vC8sVAwzqTpsqmcf59HzRPLfVPIuat3nzja2a+SGM2O1vS
bGs8iUGY2bvZMnCG48N3HlO/mp+toYr8sSt7QnT1+g9ZTXN1TwwDrR8Eb2vuI9iB
OpRezSM9cRpS0DMsbK2zqS5eBEp7xirQqmr6v94I6GkPPfyCygMdIGwDwAJ2JW5w
4jgdeEUQXyfzYXot3YGzfLFNmL0cPDJfUZixHs/JLGlUyqEjCxApI9TVzJIx5f7w
pHooqdhsLiJjeGRG0QKq/+SsaRaBMcvwalgql2sI7DvRlaoEdhAWeTPgd83bizWG
iDdMWdwPwFKH8uvxR2UiqDvK6imh/ORJ/WXdE44i2ySS2bebcYpltq9z1bphSnxa
2o/7dCLrW0GvJz6lFggzMdEPbFaG7X9lc1xy48xuFF5VuOl//qYt2gODueRm3ENW
XkJueBMa6VCI6dHWMG1tFCl/osfVqRxwyDbPNGG6M7GJho5vdUegbPY1R9y70LXi
K7h/PviSakhV2+nhXjUwDcFDP+0RxTESTzjB57Ss1FewCUsFGKecbB9jER8V84f9
B6FVJWSobMH7OojgupZsJnYD49wPNomruRw/86z7q24M3F05cNL0xdgz4+2kolW9
qP+TI5Io2lSCkNj3fxbd9muftwUD0HzGksgP0GnFDyNRX4rZ1yuf+c+h5vVYwcpo
Iw0ler0KWcoRGIKRwtMhH1vkdEEG1TxvcK1Pm7cv/b0t0exfTqSyCFX66NZrF3MV
tq/LA9g820ULwpXPIv91pSPl+5abvcg9KNGXYrpvHasbypFzUkfxp8ozmmvSLFU3
x2QmnxIbRZupQBdC3/V5hryogLV5I8Vey7XxMBCn28T8QeIP8RurD3jdtlw1H6ev
1HfcAJ9/bLoEAHf2pZ0L9pvV8PD+5nETCgCVgj8ks7he/je0/m4oKD66X/XtVnMh
HhXw1pcmNNzCv075JwiqHY/Uzv4+VmFSGz3ecCN3RTUJ8Zp2Ea6GDruipB0gnJyR
8VfTrkdszoEpA98R+I4p0j+ZJ0ry1omixwx7Omz6cy/GRxAY1zl3SHxFqctA357m
4RgGUmTmX4h+z7bnT7eHPxeeIUTdMuca13Ba/di7cx77j9vQIQaq9Qyase4LqyFM
aWTJM2qNng9yObaMIIQ/+qSWfrdmlBUhAmfOBOGPdLN50ah1rT8MGmzHwcNd3UeQ
p/C6YdyjdXa158PHZ/7Cm4ql2nw0WObm9aa1A+LkoNPOTj1oUasDqe72ZTiXF36c
oluz4dCkxbBFrwTTy2AlMZlTKdt37GztIKzTp6rwdcd4T74EdXJzwFwznOUqAWAg
RCQvhNjKms/AVwZK+zUv5GNquH9cKNm7JYC09e1kHB0h4hk4YXwcZSQ1gbbD+aBh
KNXwn40vAzzG9iLXFS1bB/B04CQ0nyDZ1KowFaKiV3O9pYLub+KEImfJGu2LfJPk
zIIrodJmlR5fXmson60eHDUdoem/LMfW8l4BcJSZyDLJSYX5EAoAKcu7VUFJfvTJ
wviygbahZbF7ywHPXfRRdD9O/YjAoWwfYpqasJwTGD+myOtL4K3btpknnS/APA5P
NQG3KYTnOkxKZrFg/cnHAcODFUfZnkLZEAXuz+VOykU2XXhlMUkU18RHqhyrxfQf
lW7aPPazAS0nSBijzxgFIi2tlKYx0n2sqgjDqwQph05+CAzbbSZEOrMbNt1udPPS
fXrSxI9pic+5C79JbC+6MuhWGnBkSuf39c/L/qz6MYRC4wQqaz/ad53OeMbi1lmn
SU5sFmirtmRXI41duj2Ux4CEBx+0kGXzXJHQN3xVRHNKGfmviNdKQ9XTM4KQtLT/
QKpINIWro5SRv4xhjK6QRZESkrGQV/SGqDcvtM8scBA1nobdcJcUKfKZ8asYBkLe
hQBljoWDQLAIlvxYA5Gb/gsVIzUbr6qn2tM6ga9To1uovyn+smVbczWqICj9Z388
UcQABK0yIRza7BEd+szEWsgEsI1F3OkG8Hwk4XQyVrScMCc6946EM/gi7/rGC/ug
btiGWUgPf9GokV2KgpUpwCQpER9oL+IbuXiUXZTuyGc+7H9FwuO1ygYW3HRpb9S3
S3jQyQNim2tN/U/entcyMvs/WVLiBFDNFNMqlXpr7i0scxYaxSLugtpROS7Cvcj5
ijZwml5muBmimxPGs8Kk6zbKiGvzAvvsCLWLx+/iJxlVySjTMmJQ4nctMcpwEOiJ
ZSP6Jtq35pTsBwcGaEj5i3/G+65lrP7y1zfjHOYdrMrI+qlxcxigSFHuzOpoUKag
V3JvMN3Yzz7vGokICESBqAxGDreZ5I7NmjkVJJahaeYz+I2YyyW+YmHjjZhdlrRU
68lhuKXKqPxnnl3YeavBRJNXhNwg/KwGDNSQAPDU/kTkvmqPJ3Btct6+ag4zd0Ve
7u1TjptOQCb2XTyyAx+seFNwiOEf784XACDH5KBGXGiK1Vxm+hhcKpcjFEGJQ29n
1wS8Hnp+d4vfNLLQhHBzMX/mvhlJmrfqVDcbkuxGYHQVmPSABwBPgXN6vUGa2mZZ
bDzBM1dDWqt0Sf+ajgjrJvkKBs+8IDhWDQqUyuOW2gVublq+koon4astEIjCCJfs
ja9wO30jqmV+bjpOEwmn+Vbg4oM3qev+zodIH6AXPEcEQesib5PIiiu6nAjqfubr
ieK0Vx79WlMHj56NMTRRAfC4nE1dp+cpW8OEqXxZdh29uO0rU9paTMDJ/OBQ6qUn
PURUGDqZ58G+SfdhT0DLIg8pR2rG1/SBAOMv6m5JWq/gaEMcXa5CsUZSjVEoGvjd
yQupAZd75R1mCnvDqN4a/tjf6MELGtapK3AJgrtDjKzictkY3gjrw5a+/cSemQF7
+GtkTZxEUwBwK/OKVyc9ICtjHgtY1fmY9CtctdiG2t6G+EcPzDdWy5RGBpAsoh9C
sxJePisqjmvhlXblE2AhG8TSBkyhZlR+kW7rGyIEl5GJ/4f+5G5GloxoCsd6GiIG
clsmkQJ9KaKbI1YiKxivYQJ/nm9xubIcxb7Tst08pRA3ZrzhyLWjzsMJWC+p/qLE
VC5h1T+oL2bpwAtIVWklgl1bN5Zf5SiVyAKXS63qSpbvUjo4JTK/lzrNpdXAXlr0
pbJHp3zSVkdDty5gRgqM23I3v1LbygiqZVzPxSSqlU/0JXL2sd9ak6cW5QLdMpHD
KqlqCPQDeeLc2nU98Py+hAZ1pP5KlrtZRat1OeBB73AstkPXbrMJTuBCwVL0qh0A
mmirsDtFnVyao5riLshcxfej2/6fHZ74HziZzF5gFSiItAGk7wzbjIzacc7MSTTX
tlhKy/rZkulnwyxub3N7yow6Biny4j8YA1OQpvkQZbL7/hfbKeibRnEV3ZF5Q9HU
F47L3dD7ktptU11XeC6wwTogiXjFrS+fK6pZqDssHlbfrhuVlhfNW8CK819iDJwk
JoXVug/ZePh0nImXeiEfBwRrJYFT+H1dVBhWzwgVWZsb8inZtD285qQXLmblkoeW
6JzUS2gjxcXOw4Rbq+xWIDD8cqZIwRcG7wiWSQwCNfddhqi5O8MWV30Ihyxtq30S
bpO5ypZ0qHL/GuySHxb5EPJ9NqubAFQMWHxjQ/4KEQqGTw8a4cm4WEponpKPCYEw
L9mWRWiKX9wg7eMoSKwkS7wu/YrADCNmJFtFMj0pvSDhPb0ShnrFnkrWdvOzNwR2
HpB361J5T4yIRblDzhraexMqaeFaPu66KsbDlag4uyCL3VmJ4fShLFzuoL4ZZzmv
CtAP+urXfaJF9w4wzuyuSuDkWeFTybl2vNebZ9yBwh5FymIp4xAzUcYrtWV9hMYk
CF3D7NNqFOj4al5I4ziUPJ7lHVyR5i6F9obX+BmkKrFgx5WJ6X8TVT5ri71Y20J0
9YDCdSVaXztmtRqW+eyasrpeGF49vQ9kolwqgyw5ydWC5lxEsFKrhP2UB5g51iN0
eAcyeXzPQmq8ScIQqSAP8PsWtPlsd2cG/YiSdKJqkvtbPECSMDEsirWZXXVEYRwv
4fATBHrH4hkJja45Hw/giuo+cXsCHaFCgB1IeqFadGnQGpAfMOj8cPmT9UwsC43L
tMK0qaMZN/5DeB47vMHdOmQrJAtxsIp/CJSRfh758vBc0eSlEGdYLEKEaxJ03dzx
QEmr0uug5TIKP9M0T6TIdP+nGPfyhzGuMM5QLaKxDi0zKbMNrVRwYPd/PzgyzrGk
q1cOYtkiH2mQvF/00CWc5jRhsajBQ8AWPvTXLp0guvq7oV0SVlub3DRU3DHo01OP
ePx4wX8WTLGQGeB2YdkOfOxl+tMQgfbaT07DfwjoK5xAxmldXeSxifkxoC0eabVl
SQAAlo3FqhMEBaswzMn84NS663ETiCh/TJSTVOo4qSAr7UnyINHoES4fV5BLuEo5
Qr8/26E81CtuyxRurVYGrrBALBEDW94dkk33WvK2Jv69u/U+p50LQsD8EcBaymXh
fiKdAME/k+YbOMnOcTTi+99eiVzJ85Q5vGlhVmlD6yyhZzuNYjman2exkfkzZhuQ
y5wZRohOScNFhLMBcXJrSok4NTDBxX2UTksBbaClJSZUSbSmCJFYJKJd933fziEg
JmIwqWGOAB47AxmMiMxyO8+qj1Xbri5eWT7eOep9iYER0HhFIxPWo55LKw6PtJMr
GgiqpNXtwhM/6kOPJCl0X81G+CaUoH5VpF+RzqimdYm7d9ejmW6eMprM1QCk47q/
C/CN12zlduvnFrQ3WeWfKtX1zgFIOOfcETCZVpFZHFHOaBPEuowA0x/cdKodqmiG
wBhqYXJkJ92kTuezGlO9h7X1zXRsJxE7E2b6/SrHdJnZ2hF6NfBDnbHLM5KR/bXj
agtKjvVkzmPV67/XijcybmaE3qojEPKXW1Zej5lOsPC+q6pzC/y95YROuSy++cyb
ArbJqJTAWDFsNc/PrtsYvqhvqVRG4O6Z+bziLUtLp5Gi7L7tnWzLxVp8RodFjXO+
hnWbhxkyeXldf2sTTKtsSkpxhk8whzEZkgymuBzIlAL4Eiv4+RtSNUzyZqIAfjD/
AzzmFjWsv7AStCFRVZgwnRD0W76MSoEnX5NPwAqRiTOCmUcuDVd0JuCu8VyHsKb+
JCwmRp1pf3jBXT0plYXWCSStRZAYBvmHWo3hi8lMvHaNa7V91m9JBFHdsxaWsHqc
cQzY80Aj2YVKxCZOUZHbU+Yvs9+i+8X4tdi7RvqA5VXDF22e8J2s8hCHxHyAMF3G
lGDOh20p20oqNzvwOaTqjPlhxSVd/+1MvTaJLaVevxQJDVtiyI+BoT+3U7eDJqzq
dG1Mao4P7kBqhLAKC5jz01nkUkEP8FbcyzAipCEbEhOOvjJaSmNDQzEoWIEUsZzd
5gWSylKfOku+Fsd6CKqBvBdG5oxYdXDv72LudPl4oPK0cG4QF9FCtKCQ6hy+Mw0t
RvbM0O3CcqM2e7rB1imzNOFXdCgQhrIlZ1RJqwIe76QyeY5y96GA3Aix+WmHcVP6
gcBzxQCg4dtgpWdKTghuz5hPubxCUZ84pk8UI2EyDr6dzoOmBbAMLLUBAjTGaoEu
J6FaH1srcwJHIg4zGBOryogge3Wj/qpEgiMhLlvMHlZe2garVH/6i72L6184/gbl
TjtwBF03hNMmC4b26D8jV1dBmM1gEj+KREsVl9N6iL2aHKdrZ3N34JblquQtrxzr
PVl8eXsd2TN9LCV+ZO0P/uONBTtL68hsLOaQtupfRMaf6Y6Kgv4QmP5VdpmodZwf
dvSyPu3pV229yoGzqFfiKMWAnZIvkBwFjmCVjJO65fKRUFR93ITIal/7Qs1P7e8Z
oWu5KE4gRzxnr+kQkcB5+JfL+uaTp8eLZpstaAL8QqLWjvNbnqv6xr5vVIC4FNfh
DGZemFMM2a6OOL1uYvimKUF0cHUNmpu4UcmIGYBqG0mVaT2Hw/oi4UvmfRRS/IhF
e+fqV23fPhgKnda3dqnNpn1AUM7aDVks0IitrkRV82T+0U7XfmGpJ0YzQG8ETAQu
SmF9i1ps4grnguAu/KZ7M8v9CMKtm+9yNVlQ8zdxSPmSpblp4tAS2E08/Qg3PEkY
LMMsfaF0BjHgV0eS9sP8d751thH2xK5xwK/eiSYO+yrMdGbl/MgQWNA1xbYwY3N9
Q2AhyeHG00dbW9kDQKJC01rweUfVAVaa3sZJiwaEUoufRuo+K5iUJeSqg3czbHBh
7exxyBx2xxy4RTP6QENxUsDBy/4R9EgyK9eJPcPMoi4rJYXX7P8UvtoV8WVOuyzL
4CvsTdfFlQ6DLdz3kYdc61VtY2eGCMvdXMPoqvSyABAPgU8WzsL5UQi086dYnNPN
FzXifYzcfQWUgnZQrQ8dRT8Wq/r3KCA+YzTPcADTOejNJJoFlR5FjFCMgpOpWCTK
kdSEW6iHU5JU4oVTIGXy8iErPfxAdQoXpq3+3rOg0t5gOVnO5f8EN2zjednzb6FV
MB/tEJyg/gHDR9zOIxzF/OBONfvAbajLhg25w6h14c8o7yway6rJ9qG9wblHeu+T
KTQ5g5he38jGfYG9qYiMcd3DmomWY3mqh+BXQgmTTzWLhFETil3igCBdKE4JnA+a
OOENAL7WPHGxd6GNIMp4UeFoQN33n+dqSaW6sYZF+z0c50QsXbskDh2AgtcxXphg
HKB91IOTo7c4sBA4pdF/AjoMAnBw92X7JJoI9cD0r8jswJlL5f6fZcfofxKfl2sR
5Q2OIQ0IrZBteprSb2rpqqWOisEy69Mpk/z2E04mldaGaPlBCvxPPxOLMdXNLBAx
+53CKbmJKxyvpb6LDIIMq+NVpJ/ERCtqZgamJ8x2N/ySKtP2AHMzqotKp2ilUpjx
CK+wWYT+txYix5CJLrBr0EpN8jGI+rN7VAGxAVfOid+uwqMH8GjW8BA4TNnblSbg
4wTa5SXSlyG8ZFDslhBTZA5bq6G0R1XbqLXLBDeDIJODPeXbwYYCtAEqWbUneq2p
SILFCl0n/HrFb0URirGmdtf28jQRTpCUFbl3/e2ku3ujNwwxpnuAqKuUleeMDCEL
cDo+/Tj5wxOlwymODOftWnv3ze7jp1Jc9pb/SGjRqwAMO7i1iyrbYCrst3t4TRqg
W3XxguffJe+NOo06wu4ED36UbXqT+GMi1NLO7jbNCGGkdrNRfC6r+bff+5GZBkdm
Fv6ws+Ibn0svUOM/CJ+QLA9B50NSrqX+yoadx0Gsp7LoR5Nq8tWW1Cko4F9umHV6
5rUXeNhL5dMFtuvexetjzT41vSBtIeDD2FSWUri+nS0KupmdjyVOOMKxcYXCLLsk
THpRrAr/0nZIjrAzTFrnbURA4oO75to0uxWM2UebI7NrQQPU6sSqKG1NWPF1I+5+
9ZUSNmGHrx5LTRovctRp6QOI/bOqJOpEoML1LPbN7oJ9CA/P8k8sL9kgljjOSQlN
PeHj21Oe41kaHVU06QZhNrPRNArA3opZl/ruWNsohB2/58CFCu1QEbdcyxpPraHO
ufAgv298jAIM6lY6hhFuxipijKlIz5Zc3LyG5QESRRnNSRmADWESQzGctL4/SdWk
M0w4w5jgA1m3uC7x2Bk+pURlsaPTFK6ycg4R6+9Pwis5hp5Nd3gwoCP4MF/KvlLm
x8OAJJhH2Nycq/+2gCv6gVCIjFZyxXGB7S6vHHKYgwdx5CzzkEh0+VFKET2L0Tvy
dP0dt4GRUglz5bJHdupY+pSu92rn9T94N5fw0v79oMDKP8cXTEyf/cypFfQ2BEcv
ccD1yhOXZUt1BzY5TxzHsoSAeM+GVC9/nJbWA16fPBN9fzh5PPSf5qzcqa0jm46F
8Jg6GhnoHdcjawl1WQKB2JQz0ca3b32TJ788G089J6rWdBeqfFxGD3SS87H5Unsk
bjJxfPLDj0y8VSzaw72V5lWxsQGOpV2PGpb1GX9iVZ0xwf78Swkq2vTXoNxgHFqD
5wUHhanAWhQCqzYqZonRwCaqw0en2yOdOmbYHpUPu8+T1oKgA6wgIv6D659YCKxv
1BevBxhlmBQJKocaUmtxZvvgsf8t8GR2FiKS13fhbm9MUyfJWvBhE6oWofrEE6Ko
C1wWHgH6bX6Ea7Q2ssVB7Ilxr0RFqwC1exU3BBzHR9RZcpH3GExrZ+8hvQKeAvq4
MgOs1nm77LG8GURe4nhb3gTEolIjkR305LmeXEg2zb0UYXouGeuQ+z0PdczBTTbF
+ZiaX8Qnn/VW9C7SNNRPvOz11QRW2txto5o02QgDKzshVX140369LYz0K4h0jS8M
EStR1FgG5gKP9R49SPIX69WFc16L71rw9PoUslqS7bhGP6ANWz3hLNY9hzzBiuKc
T8S3BV3AAWKDpC+lB9hNu1djcuzRsdIRqLgks2BRxK1FhD3kWaOo17yAPN/neXuU
VojSo3usZrTkk6b/8kkyJdxx/mUNGT2yyl92KBSIcszNnSA0m5z9XfdqJRBunx6V
34AwOwrF8YHHfERluDpkwJlTJlQEcOw9E/+cZ3g/RjfR82qfLLakusQ41DtUS9CH
qjF9cFLsA0iVUYOScpV3/78IbaueG7BWlsWyfbv9C5pIb68njR2S0IhlmZfhR0kc
JrQsJElhq/0M+qhtTR5Bu9UQ7JjI9/ra0HaPYZG5orQ9E8pSAOeel0vb0noa67bg
pFFe+eRVqRQSSk9OGvkCXGpUBhhTCC2zbrb9Ubx+J/8MHjON8xTDdApc1CIuaqK6
AIJhceWZp8FCuYdD+dL71AYNSC7a3opvFh0Tk/kQUMCCtF5Zm4sLGfEiXY6Dr9bP
KhK6KN4zgInOJLrYmSwQbD0SyBsvrxurT9WTEQnThntIz/X5Qrt8xsHr0PHUxa3T
TXOkSYWDau3vhvQgQ7dJMzwQhUBiyn0Ul1DubWvq22TLPt+rxTmvMn/XmiQc7DTE
HfwDn6AtxRpPZxvo1SlkJ/E6yxje5Rgc0yqeIVt11FnzhTjZ9Mte2fBEkJzvH+iN
oPbBta6Y1bVTUPLrCNKX2S5yfBBvx6MQ2/UF4cvUqtVxNuSAviqGlUs4pU8m5wUx
llZNci0ZrbxmkJgfz+th0EjesgKhk1EgvpqeTBqfKZ5eqNa33QJX2X7df2bljqD2
A7w7XSUw21JqdR6IrD+WYwhxdvj7juMqi7u7c0P8C4XSmtOzZj/fFDnVSuAPqWJ7
KRRzUI5HzDcvj8aDcnyPytTtUp1JEgTfS/nY1s0RylYkjT6WtAL1T2K53tQMKwAH
KdpLRnKyNhi3rc6l1Auk2hx9OnGh/PGoLk1npwqLHYdSbRtebhYXkDL/udqIj1NP
7O8DRj2B1kDmft4MKz4+yjxFFWRNvT8a07Jx/fVSBTdUo3VWmvhekW6w01jTsNn5
O61pEvoVqW2gvLNPO4RTW8xU89CrNWBoYAKUG8ecxspE2phOfr8yxLiW3GWoyZJF
ouO5zSfOI63VrtSBUQ7MUKuYY/plKUap6G3Cgs+EefNpGB+qx4rZuVp/6RLbTikG
DXFwDQGClFdWxkX6nQLGmshAnRAsE6nD5baekIA9e7Lj1OR2nxhpr6qOxqRaTdR6
vz3TY3zcPIdKdfl5pKEGJbWoI1raszjsLV81xia2Rh+ySEnzTmOw9fuWJwlZC5Ki
Yw0b24IjpQtxl5V/JIDBcvzGjWCJIqc8eoDe21t0a39bPsZBKAaowGvL+I9cBFqU
WO9eFarJIy+DELxH0ytjoIuasmT4fCQ7sB2MeXlurPEqHyfVSC/eRgFtFNc0BSlR
FwKZZhK+7D/EaYEKZhpZeialHo1docGCcITuQ3LSN/tmoygy35Vps7gIqmxSjbSt
8dgEcbInYqhFAQxNHwtV54izLGByLDHMvQVX9MyXeZZYlauI0x4wfVQpXceATgTn
FnZLCmYzPZ2GiZV+QMXkTltaJ3tuhZb2babZ9kC7n5MER2hzZeK/noYLn7yB1+Ea
cCcWgU7NMOmXyb9wm2tBdqjzyvnpg3LY6j6Crm8h5esUYCcMKDsZaiI8/fgReAWY
o3f05AaxMe3w5OggkHZhhTKgvSqX5MADbz55frQuA8sjht/GqwCYlouZ834VasXX
NuSzUVoq2+ikhUrLybOKiVi3bLqvRGaG8arGblTf9vOF1JvDOUJxCbCjz3mMLLCe
Ql/N8ftg5RNTJsPwleiQ3u5VXmlYejEYAwOAivxRNwrxiEjhtJpJg1jyD30muCUZ
gscCa8Gz4uOyqFU2RgOaVoORKx5DVj6ozjxbJHVDY9YYqczUygTBvEKEejQrPKQF
bxqX9o0xpnJ7D/jO7M4478gKUkOT5pq98CEIw6qH/cna4IBvNl1KqGSbBjFd3Y6L
aZQ8o1LYUwYISG+0HUOuk+1Qh3VIxltk9UK+XV8qSMJTVNEIOM3+xSC2ce3+36kF
JHQPECC9jFcafAFfzOLhuO6oSoynekCMLr3NG9EPGUAMSHuWf9YpkLJs4J7GTeHe
JFFuCG/b8nrRfiVLq5RhGBe0zKgYvr71WYaY+wFobjonPLjo6nW8qBEjPJAKNhsh
haFY2bLPz5lx4OLPPRatszAWq816KANHr8eXYoU5srHBeOq1zgqM6hACJ/msyVlg
Igqu2juoIyaVQ3Y2tIFLuhdMpZ5iPUr0RC2B06sDBYXLpJmmSb5dG//b3BuvA642
IrMzVbVIyYJhEy59EjjEKiTVKL0ZchGL5nvTkPOMf+GjG3BTX7Fl9vIjmBlN7A/R
CrH8AMWSrKmHme51DBnxXlFWI0FLxdXxqFt7MoN7C+YelcUplycVgTtR2JRwdLhw
tO9QlldxDza3nycM2/P8bb0EUf2ro045qHrLJZ0A/B1+m7oiYxtJfz51rt7TD90P
sJl2hnWCSr7PnCNHzMU2SwHbq+eIfHfV/dtxMcnYX/0wg+2GSBOYl34wFZpaqbFh
c93kBRBICT8i8X6n06ym3+QbbhaDivwPaAm/9qaJxuNoSfYDvnGTjEr9P5+WPWjs
SA4b6v1m0qKdr2/UzMD1c27GZ6CAAc/dLT5iibvgDaryfy/iqMzcgoxZ+o6ughQ/
TZ7Y0/PqPXKlNqKaftglnxFiW89QJHk8GQrsf43YDlFbR6dvQCHft0GKaQoKlq6O
7c0vT9LUM8/o9+9ijJu4qcohB2YKZIZXg4i2nBn3tJMYRUXkqT4RNUopG4PTMZW3
la/GJfsVaMEKZiEIiQTfm+QBUvrQfErc3XwkWki//vUlaom4fHkCjyJGi7kRhrEp
Aw63btcWdKYGasu3QNQtCb2hoLRAUL0rDaNNbFtfakbD8GDpsrGQ2Drl7QhKGXyn
Cgj19U29VdPx5VqrpkbjGZm3WjSFPOWeMUa4Vn4Q/zRIx4obRa5Trsh2fZIwcqA+
QGHhCazepD7NAZXkICkxtLyAvcXWs3RafVyzPBk0NCodbtmORHaYXS9Z/jeXsktl
wKbFpgqBFWokZ7uHxjhqwfE9eLoKNwh8mG0hBXa/EBL/FIFCY8pmfHixB/HQV+FB
ogx+prhHR3YdGFx8EzRZZ5wOiUnZpvMge4h18OfPZVCsR5HimPcTPueZNE0E75S7
b+3Wjq6r1DMYXRirilEDzBOfRV10Unpewv0YU8y6cNrIeg2SA++dGJNB4LevW9rY
QBAf1hsQCv//ZaqAraTR9wS0lQwr7GSIFnkGWzsSqSNZgDRRyp0L2Mo9A8fWyxCh
zRBJiYRTFFV3ddEIqMlPltumCc7DmXwnJw659/8nEiZ0yDPvZyw9X1lkbIYwy9DK
5BToHPGyiHxH6OdoaMHX8866ifaU1XBzm6WNLpgBH8dr0q/XkLKFr5UCWUjRl8a2
FchDMzGJTRvHvtJdlw21uy0Tg7h6QMHiifvWvFwoRZRK8eHui5vU1DTswWfSSgKh
RzBv+aOTsLww6NTkOhmABrPvC5M7ZDKeyl7JH2dqtfBsQioxJXsPFk3udalV7qqO
u2B4134rWR3tjLOceX+y0fs3/2FpJ84qlcFp7/7UzkNiV8YdmPL7PaTPDsv/ocmh
GQU9fhFDen+eXkhddN5GjukkSruSItqx1A2fenEUGBZ4T/tuF9UllZvmMwntOmMp
0Uyt4e9BMjZ0S9PkzdvAA9eNT2a/Cags/08CO/U1RB9yODKscw2yLeFLZ72i4jTn
hMbsZqt2q5MtLRkt17TVZ/EetCmxnqPHhzLt7n57fPI+WsSbXez5ffCDEUQPmDde
/Epi1J5AuatMQco5Byg9vlCsRYUsVQAogZZKt6X2AWNLZ0fu8xZHq228/HCtrF1C
s3xbbpRcg33xCIfcQc09E+JUoI2mKYwGppU0h/g5q22Ld3/4gEUHo1PwAedliE0t
+wgiZ7RCqI8bSaLg3u6nGQBvkyDRUw+rV3tVJDkia+SHiTJuOBeJH9QtQEd9Cc+f
IgTX3TcbLIgMAwUOxXEobW9W9mYeWntbj+gcJwZ6JJBpqySk/cLWPq7XQPwhvC8v
gfilCx59Pixh33mGW4m+xI+jrCYVJhWsAoP1qamLydtfBdM/3NatfpwELmjPj4oo
LXAnXvvM30meXclwycBdwwTyuGnbj/+PdhEvN16Kx0en0+Q0FWZkIUFye3aIuf/Y
4a0iNCZvuXp/9Uf8qfPMWSZsRo6/4a+TsTK0Y94Q02pgmV30FLsMcia0M0r8bbGV
5SmKr5AGl0lWx+rTecbzeJCWVbaZPp3n5pkMz4q3CRzy5eD2JZ80YPY0SFy7k1l5
holeFmCmUg5PgEeIaChK5oc/Ln6qn/+MIMKCEU7CeB/KdWGv2waPrnOtCLSjZC0k
GfU8R0pZgQ7oZMUHlsQS30J7G+MQYAEYiMbeOzslM/v0vUBo+4EYqtSyaIx9Yspo
lqwislthQQz6xu5UOYv3julQg3Kd5H5ikCgk4vPmbSwZnTT2XwhoE8K5MwXkxYIS
6EPklwF/V6fPkpr9kZDvddr5bh605MrkJ0RxiOWgplaB/kHhwpN7gYpE5b9Q0/Xy
gI58URRxgE41egMVSlgz/4T3jCSX4hXFuSiA4Kq7sakTaADVdOfDUV20zNfRn/5e
8F2uJsh6BSz144RUme5sLBPkQfk2Hb+GdSBFxyUNIeEWgJUTEA/3W6/RPdSrZBa6
egqBg2o/ya439af9eso16C0MMOhwIa7UYQ+YY/qjpeXBBSaFqpjbvmsfPoXIjopC
8O7bg+1jkMKygSfweYQICQWeREYOuL3H7DM1OTYvrQypkStSKA3UE+fipeJ7wj8K
PV7tluRRIw1+BFoDKn1+3eIJQWwacEt84dfjgfT3QstAKVxVErMxeyCqueJMvvL9
bjeP/qXe7kwet+J62PjdLJnEHIzKtzEC6OrvRfJZXgAvPo21dXUL1SqrNMWWCovr
mEJcVSOY64F4Pvs84sg0a9DHkJ1v4mH1e+UktIZIm7+9GDDirJlf5hxFijEEiTEw
NGB9vke/Os3282DAlXUrRMvSqJhSEGv5izRBCJc6Dlc7MdQOrRm3R3OZ+VRYzDcP
gFvyWmMeqKoZ16Ri79XTueNEcEMEKsUJjpdsdKWAP7Wn2714j9zAnVvPGheYc++s
IOS1CUH3tgCj8H0/3zNFEJOIIoMo4g6u36HKqY9/Hb6pOcFSWXlh9oNC3mnAoB37
keae3xTx1kQO2EJdi32jZJw9TUnQBNnloa4j3QYyvWrbC+D6qM1IJN2j6EC4rRC1
oS2Uu67bu6r96k0qCu/HQR+uPpL3ggXyCOdKX6hnMXuyeWg0DUQld7Ha8XzFKvLo
RGoHkmiP2Qf45tMD3t7uQIVVEhE7/niyEu35CPtBge6fFG8r13kEb+ER4SybwyG9
UAscMsHrwzL1JE6ZRB6jaoRQ4aBDpHeNfVH6QRGP25UfeOCSwFoiZbdChDyuHmO2
M5Av6LsGimdlxgW1ya8iJdCb2ET3yNsxl/EfdfrUkC4VP2NxX8WxNTrWss9TCaZZ
XfwOJ4qRj8a5Etw2bp86fJtWs1NWex4+SB6FTn9JV534X/pT/+6FXdNg6gHcVN3V
vk8896QMXXXiegp55Dm119RYadFYevFFxbHQ6wlls4+L6AOv+kYoUKOqYpJ0halS
RS6AmQJeIgEGSUnOQOTYBpXqDslUBbw5WTXj4fVxwLMBttQLyM4wddi5duRXMH8F
r8LtZDIK8vhX5xn0xXuGk2A4trSxoMkKniaFXDD6d/zYcQVC952WWWttPSrODEav
xCZjD1OUoupkAP0dDvwDmX2F9gh1AqRy7FU4aW9opgKAhsmBTPPxuEI+ADbtpgms
g7yYhvZVqcvnkIwi4HyklrIoszHPSalzNrXJ8Ck6zpFxrnFCVJIc1AKushz/3J/0
uafIxASSOovWvSasSHLp4cNtTPNmsOlgn8WwBmSQcwnotV/cj3LyN4XfIrkcAzsr
hSoWujchBCBKKaPJDi7WmBp8I5SsDlAFTsccU/cYER3oafftZpB5GhCUweYxxsch
b6X/YAuCJi1Uc+ZMwN+zlz+P67lK0YGQnXQ9en6MMgqlnYATiXaTH8R8GboMUiLQ
0UFT0EEKRT/c4a2bFRMjFgTA/6lclCMgdfAonWgZnACO8CifzsVGDdaOcAYCA1ou
meJx++RbY642r4d/7HiximarBgdnnEQEE3frtD3GJ/NacnfHWMZi1VSHI2r/uKjA
lfzBGFt5FVBOe97JoJoGjF/Ef5I8TyQ24CVVSbhhMyeGq+/+YZ4G4ZbTvNHZxXM5
zrdzeoYBuVPIO5MW9mLRybz8KNybthhLEsiasxiDMBwgy84lPWTCSEWQajAOoRjz
DUnxliGbcnQfBQAENd+axtU0ndXYa6j/5Afj934o1vPq9mqj9X1mLUouo0BcSoO4
1pSqayCiROKJKv9k6sA0ZfcqgJuS432d8P+M2eOD1rDhwE2X/yCq2fTNDw07pnKr
cnq0iEIGufHgk1oRdqt01pLCD2Sm+qFha8GHi5PJLUTvaX0YdiZpqqRDCb+canje
+ixHhmZ/jBjGKREHbG9I8GMGQwfZ96ssOPuqLAyZ5fxZfzZKOlJiw92ZYvBqEboS
OyNgIXywUDteyt5gjGr1J68xC3fqMMy+6pLZwheNKDXAr4Rzcm/3/66vNwK49y5A
8cDEBix4QO4XnkBaAG+fXkTUkgj/Of+ohVo2YaJd54B/OWd/Ura2Xe614ddv4cA/
1RpB+x3U+Hu25HKyKAni4XctZY6VN7ygI8bQ14hsti4va+THBy0y4oRBEJTWNSL+
J/DMMpOmjpXGt2RWuQf+Af2WZKYOP2LsCpDIPwg9lq22s+hcTgp9DfOxxeFVcN0D
H0/9pwbHlaIXImQerS+GnKa8US1zZD5BqnhKBMpU8WbBSmPpLIon+0hVpnIjIg4q
lG+1lDn/DC5ji/5jzhSSG9EZkasM8YYfRGU3fYDjA9J5shegNcQDpmFlTaDqeDhF
jMnwEpYLIU+F4truucx0M7dy88NX/DxFB4ejnPqgiJQ5VcwgbWDp/LHTTDRrUrO+
Vg9ccXaRsYBR2Rpu+ljEKphzPlbBh491VZWwamLby4TKSv2WEDUb2LCJyrn15e4Q
nPdtQLYYuG9mvaY0MPRlZ5rQILlE0epBPgIosm3SoTWT4cEq8moQTO1UrYiPSyGR
6e5Orl/0AaCUJQ6FWx87HYgYXCRbuTcJ82vAadDIbYib3sMkTnhWaTFEv1ETknJR
bT5FoK8e6ISebMVxFfKCx8eRewimQnZt2qXHsKulMLJWbT5oYPaAiZyx2h7GIklP
UCgREMfGxtxHB6zmBzHcS/w4X78NkpgO2f/eLdRwPRoBujAJuKsff3BdEnaopIBw
FQ4s0ZHOWPYcf6/pJYvficYs5VduAhGofWFxqcodwauta3rf8jTOwERuknUa2rHV
VpFJoX+jbLyQhVmnz9uZzpFRlSfVsGypTqHxpjVzCqyioiYKslfyPD+cNDEVozKC
aCClSOte9Ns4zS9YSVwhDGhqzPmEHWwqNgTNeKd/LDVOqGtpWT+iOX/A9MZ+XS07
z/ZRI9KF4a9TQ469qmeTCoiu3unuOcbLJoe+ySdd8dn2zU1bz4sndXHGYueUciqy
H2sc9I6h1BBI9Z1P1o18e/YFow5EYGvCUG9HJrOunrwhgxRMibKG4AsvnQxNecTp
iOEJMklTxqQjyrdwKKd4CsTGcbiWRQpDKTrWH4VNXVmpIGFiSJVg0ogGSQ32ag6E
6Bll2TtaLwRAZCnTfTG282Kz47cAUoaeuD1Rhp2W1oFFF2tgUAMqWvEk3q7OxPvB
5Racj+r0A373lmOD+/sxK48CQZA40yYrc0Eo7rFKPEMvNA58XDtC3915sUqvuiRa
ME6hLtkwzJwprQLZ6vvV87LI5eDxW7XIcfptkOgSBUWWWhv73nMRblF2DFuceV0B
m2JgD8kgwViL+cdoNaj/18dD1X57oCxcp4S9tWHqullGFF1UB82XG9z1vZhFlPga
LOV/SVI4yxHNJN5QWQNdpW9jRhrq+t/KUE6plZhERlN5Me7aL5h3SAU4ZOIyiqO1
2yX1X7Q09Fq6dncUxaY8B7vcklFJta8R08ETJX0qc55aslsEFYdAC92C99/Vy97J
uKaXHmzrrFSQOjrQRytfGp8HvwtiYoa+PT8r+FFpu4PYNVNDgnYiRFzENpWPqNFN
4tnINLpdCDMq7hm1Z0jS/KHUABXUEXoHI4boDX7yHgwi/jeNRKZAOvAVm+Ncycpg
Fkuj+KuBM9MVxLf0nVwgDHS9Ya489ntXuaXzROWAxdUkcqrPpi4elj/KPuKdJ9a9
H5gN6BG5RY6jN1tJ+bscJV/u/tMEaXtT6BH1mRaKyk4NpuPcZPPB0/QJnecVwexV
KZl4CkcCvdR0mzueWhPMFY5nyn3usPYym9Ua9SYCPX4hisiW4Ii2YADLhoQP+AMg
vW/LdXyUEli/tY7nM6B211s1RdLxd38Xfd4uyXQd4znVVJyExsXeprtt8ngVUmqN
DUMHc1qRBDObH9X6oO8/Cn8/vKqx/ioAjm6bssr0ag/w2Suk8zG0v49Ra0bTLaqX
0CTLbtYGdal/HTTvXO6qNcTSDkLBEyH7HQGJZTCJCBo1IRUHEpwXou0SsCCY24tV
jtKdJtPeJSE8zyyeTEf6qn+6dGSv/exJiQndJYXwi9WO1kyLXZUvBpb20lOPQzQy
MgS+0j+9R8iyBFI2oOEy7tgFLLtQoB9EOU5JzSRWZWAF2BEfLkyje0+WL1IBd+Zo
aKMTPIroL5wsjSOlGgOUkZsyEIf3ZrVNdhnT+wSJXNHHSdqiEl+Bn9norjJn1nuz
eRSibDeZVWhy0h8vTH2G3MmFXX0RAxXwQsEzQahZjaDsXXRIfRqav+3CoEyNdbQP
2lOwf8mSiu5iQd018tUaKJlZM9SNDj6/URN7OswKWYgaumhvrBpLh8NvpviOV/5e
NoC4AqU3HcWhy7sC/G1WTAsJH6kP7kmg9mffjpfoxz3u7B6hmfootdeEkKIA5wyD
XR/mUJkco2bCT+M6wITPWlxHGbbU13f0CSYd1O+sF++vWunNTR/vDK4oaXheLSLz
jPq44L9JyOVenXAXsXBEzrYFKAyueiImp0IElb6jD3ReHvqqow5VwWBByqGgnOQv
0WNJ9ptp46pBx1EZT1EHLKN5p39lqCB0fsfwYZw3/z+jNUvFO/aGFeL8HNBXVb/8
5N7UPUCJ0SsWW6Eoh9TyGob7gzFu4hX3j9LV7ULLfSKL3XayXeC61lNX4hDPrlGU
cMaU61/39MXed66bMJ/vQfiDP/n6gErlPSWJYUwj5XHkS37nLPaHbAF4IieIRo3Q
PVdB6lLHU3onAXju+Dwst4c04/9zBBIH7BN/JlO/GrHvl7Cw4ZTsxyL5xYg1M4eH
GA0G4su2q4Zi0Z0j42p0C7iNm9JDhS6LqiO0lVxH/moeHSe49ZpnKlnPySvuHNdn
MZuhei7JW8ffANKRsI17qBb9G4xIgljlTjbfZLsx5dq12SoUa7a5Ct0wzvONBuPN
LZU1NXqO8Hvw5kckZen/dQqpUL/N3zhn/wxkNDKv4jila8kVaPtp/mbST0n/vf8P
Mja5tQU5VZJ4TSgTr7CL90Q+ZYzuvW9EmH4kbRzMNca7UhDNCNeyQcOBXn19mTmc
Xt5b5YEbs+kQALgO/JM2boZutk/WDzIrKIuvyEM/epW9+skTx1L10EPEMh/anYbT
5nlV5JuC41a7/PSJAhI9sLtwQzXxIAPwO3Ytpg8ajyn3wtF7oi0v/8Uf4nktXy6e
y03dDKaSgEOMX74htLrvlKlv8z9sb4B3L1uS9bhwg6DOWroX3HLHqTWz/hn2SnZC
/RZoO2FkbrPaXHjOGZ72e2zSDUkjwJhxy4A4VTOtsBhZG8/sKUMtS/E5KIfIgTyE
LZOjwzMsQOyCUWrPU9ulk0K3xK7k6d8mzsNmss6dm7QGVtyIdw9LASyHwObWdUJh
n6XDbLCOvWMugREbWPwcPkoxtPdet0ynAHxXjgwXu4O8ZJbPs0Lf5AX5yfv2v+w9
o8JI999I8L7qArXYXAtpiq6xfWDMsN3lEQlor8P2JoXWYBL9KJchSnQ2gX5qa5Ji
JrJ/gvwytmTYaTz83IUaQ7DV76uPTzrNomboVZrREbSE38/wABuQHHSxjUSUsjpi
0fMv4gHBdajWwkS7Gp/KqKKcDShhpsD2C88v9cwCVYiOAWyPlPNLaG8+dkjbUYa8
tT/LzFwF8toFtnw8uJw2gI1lmdxYWB18wUeGMu8WjkGMc6JFklC/hPNAtu75Rth5
BxRO3EKUUVeK1a18GS96K/bdBbtbBqmKUvILmDAdVxUZO2HVbZp3AhJS7lfnUho3
1gAVObTwal/q2+DkCRu34/8BgzlBXlHXKYiaDlNl3X3WXsI7x8DxnBvn9syuhs3u
szdpku0y/j7g67404WfIc01MIT4iQMic9oVt/B1HawrHe3uyEidq2/H2EZxuhLfo
UQ4mpnwPHk91Jtvdd7mFicihSlPl/NiH2hALRcVT5ZvjxJeJd/XmASqLOmMiRpPl
olxBPP0slMqEgHFzY0HtZHbrmyG5uIf8Qou2PvE0Ej/vvet2TzdR8NR6hnI0VKwD
SJFVEoxbGUDjPYn47Rafv4vWweF4VZI3HhzZEeqYKynizn+EWcA4iI5Gv6kIxl0D
Ql0wJGn51xP5RgYZ/jIKC3gK3zmLYmnXex7RRxKzBXis4TCvTE4GQBaQQRkVUgpq
5XLcSnBLTfLS5gboPUdNR9SRd6CqwJofCQ+jWEpsNeMErAWyUVjP0hA2FwWKIu04
b/NIXJzw3r7xDBITrYGx7yDFK89mMN5hCC7kUTF76nmTpUZ6Jjj/z37ePOlLdKs5
9HhYemo3iwrirk3IL3Esb/ysEAJtSDC3VvwILOmfHuSpoCkzYSMkvth6Lz3S8YWx
+KIwEsiYRAu6YzzIirpP7ZXl6iOQp6W0OPKnIpC2quv+IN6bqbKW72lzF5NADTCb
mWXBOGXNH9SWL6HisVmNRSGNNwe2FfCa/1IaYNG6x68BuA7w87eva5rw5FEK9wvY
mRZKk/4PZY/Ez769PKTk1665xum9M3/11iFMhwJURPC+f6Q9UUv3ho4k1z8v+ILQ
HOsH/z9AkIbBoAogdgE2VklXXIEZOLdDHdmyPCMFXV7CgEfynUKbi1KPq/JJj/ci
cVElv1KGpqA1ZAFHT8plXYyhDH/aO38lST6EtWzkECF75Z7YG3ne60V+J0KZvQHV
88VOYZiEnUVoBNQ68MqU+6bahYA39drSMp2sqSqwKXQ5WTLc7uX/is9azbpEYdJX
mfXE4CySmu777Npw7bP893Fs7OWeGUFCsoodhmxUN345EKhBqtFVIjIncqQvtAiZ
WLh4VTl7RmqmIJa3LK31D/hExj8HkFCRLdwmsV6lD3NAkV1JslHO4YJJiFLyR65N
4KJPr4ZcYeq9l9lpM5DqJUxvKJpCNliC/Ye/rfk5/4KWouA6aNeaXxMQIypwWFLS
LZjfgANp4O373T9VVMMS5zjaWjaDxo2fqLP99OO/aivnY3KEV/dvI+dARWJOxEx+
uFeod5iL6Sc5gdPPlHu+UXytSI+uZsA+wN8Mmi5dIXaASPx8sdjxMKeDoYIBAeet
2JwBxdzRwKMk50j9+PXeuJjLwQxEJ0YoEKYcMuJZEr/PNFjq5TmKnxG4ANXq7NPf
pB91Ji1PGMEniGNYXRlI13rz1CDvJ7Ee1/ShWrnmUgiK/UqgDFmmvzUakzwn+3+i
pi0RI4a9/lvmJBYg1/9AWiG7Q+YMNKx/VvFZA12dilVg7ci+2podkzkAjMd8estQ
+kO72187QICSvZDz5Ew8m31ngXPeK9rV0GWVgDjxnuNvsO+Uq8sysBz33dcRyxHR
PA/N/L2YjwyLaG+bzpOyoJScEpvvT9JXQlkxNLM1plr+kdKZKOyWC1O6c2wGJVbW
STAsA56gHE9EDqrlHJFqIVyu2bXlJakExDufAiem0Fn7L/xO8d07CwEucu5BEUHe
wdAmEjAHS9EpCG0cRuxBeLbOaYOfWOJ3tzDXfG4/+/mbLC8rgtydrOp6YxtQWlDo
EmwmNrMHeK3A3Aj8RpuKDKNf7RcMBJcDYEqM1ow9cSRwRBqQh2K2flNrSZIGN4tv
JN1zFknWDphI1PPJRjnj0dEEnsc2vFm3rucSzTUoRcts7HdbSVgUK57y38B7UXAl
7hwGT+Uvcma4XR0HZxdB8tC7agZimHxCR3jiU+gVAa35cmIqx5bMIzDCHxBo2ZMP
E6muvUKqwrdLLAVKhJOdmR5PtokGoLHqYBpUARfz7xVA7DLmMzUrQqM5T6TXbwRJ
3qPEciWU+mKoAkJZzkbzy0F5eONAluuyDWwg5HgFqE2mXZy/vVeuzaIY7wA3vnVJ
bbbSjCH51PvHvXbRPTtT0hcGuydZmSweh0uE0G6h4r17SZeJF1bYzZowszN6O1ze
jTkHjoMBRyuVf9emLjQlwlo7RBDj0ttksWgOX16vnTC0WGzOLjZzE0GAm43Q801j
BdVWe4iOOOktMw0LVMEphZgcFh7Nr5ASiu8HuCkEYUhBLQsEdYNfoi+dpWa5LZgV
tXRrWvuSgjhgRCHmZrvv7FdWUHqYHpQu3ELU45yzs5L2AOZTqN2evMcNiOHPX2+S
UIsmadPrDAzhPB7xavOawNhviwQJimXFD5+z+pvVtu7WCr8DntQLCFXqbACqu5hY
LiableaqkNyTy4YkFVZnCr1NqvbCY7GsV57pml+c77Fyh1BeubaC7GXKpo3iuSYf
J7NKRWSyy84wZ1mBrnKGmS8zyrbT1flheldKSqzbZ0/CfjDHPBJvwddNuqJ9+SKU
c2Wh8hkOiu48B9/uDfJUwG5Xb9RFNGLjL0YUyrS+liknU8Iy8Ld4OaJjKZ8wDLgo
WuIFt1vor4OT14MY4Qf2nZtj6NBpNYH33vfkjS8L532arBH7Ua+bYvek6yx4sC2j
6uJ7Nv1A4Ek12+aow+Uo70uTQ5XmhzxAuIYxuXfjg5mdXu3GvPt0maQiNW7ylLng
eSmvWARQ2zuIlXkNdwEJ6rcGnkAX8FYXkqt7FoTpFH00jd/aI46g+XXJCi7hhdY8
VBTAkBU5BOf46+2sLYCsBkZ1Jrtd5lbdll6LY/G7d+gA8Tf/F8zkqlhcIKmhobGb
CMH74a8zyOXw/ZO4UyIpS6HKPBaSdmhvyQ29SIQQc/1yb+fYYy2bKF+11WCtWtrM
TVPVmfAZG9VXUz645pjOxIjh1pCNwBPLn8FOhL8avVdYjsNzZrqFa8UzvfiaA7Oh
xc29WSFQ9uXfOJC/LCzwWWjB8MQTvxdDsVcmyxTGVwkY33x+vqrh3x3coZX6ek69
cxU7ZHsqjD+0HrKzvKJxTKlbPQZIhnO9xgVBp5o8hqhkKWJjj2jbcBi1UzPjDn2X
aquxGfY3/evHOqIPPfQw5dZyqNFVBCG3Yh/JOikDPnt+4V3JlmtWQqo4aYcNKkAZ
0ahC3wk5RPEhyaVudzGC+OyyMhtgSnta8qIPLiEIAXKiBUBA0CjSw+r2Ns43W+WY
+noOIaCDv5PC+yRMrmKv1tuqMfRD6eLf9Zcq4Ikd9cFlKTmb+04U4yJwkr0rZz/S
UG9vo2KCoBsgv5w6srqZ2o9fulnl1BTDLqv5EoRPdvbQ3Ss72hwPLqNf04UTONj8
3MIriuA1Y8W+ZiseNpUQbTcaqvrQrQjFUI2I6AKNWXZrcrl3dQC7P20NbbANdlYg
4pKroW5QbYr3LT4E/UaRYtD2q9js6ETUenukOrF6vZejA/yEW6/ORBDVtHVFpzKL
5ZpioATCw3i0dPCTuA/rIf5BrxRvv8+nmxKKvdkujj0kaD7IBh44rumVH9a2KTeH
3ZL1bBvmeaK95gidDHx0ZJyelOj+ACYYUyEPaqW5nDTtoLAyqMAJJId3+LsEMxUp
HbesYeDRHV3J/547OMJ4JX9SgzGpewQSsa8CHHDrkra7gSjDFXi6mx1Vr7I/+lyJ
3AHs2KOq0v9BSBvnvClvyBw9AH4jqeGWt5mazrc6+zWusf/8pi2OzwetHzEaoLFx
sQuomWW80pzJ/mXIeer0QXvCQE+Z5J2NpCudCzTuR8hpjcDKJmdEtkSHJu7NYcQw
jvjMSrTRwEpj8dRwmDEdPjThzop6Y6AxdOHOYrnty5O243nys+jlto+es5RJ0Pdi
CspwJEqxGb4eJYEH5sXvEKpbL8vAwl7sfgHUnA5fsssb4hHJVoLumKOvzRJvlby6
/M3h0HPvm4g3gTrMmIfarmrFBq5nZ24iVQZcxni6PeOkuqCIAypvbyFVj+jg+/hk
mmPJFsLNDL9nSd6H8B56CBThcc5m83KB37NpCV0tDAGk6T19Elf2m+8KTNhxnjO5
ER9Vg6q2afXiUsIKqSw9qqM1w+iCKAruBbiJQq9jks/2eIYkab8jQak4ps8qGCKq
6j2er8ZJrYGiRL4rRr/tCupl+7Bh8V+slVmRolp4zeRw4tJ5olkx9cTuwpK5IIXD
fE1BmxiyXea1UGJzRY5yiUkl9RUmOMrh/jPxvMQovz37tk5fELYm+RBE9bt6qchB
6FEiuDY8i1CDhAhiea61Hdkzd4yXgYaLusTQ8LqceiWLuHaluu09sfV32Y7JdZXw
zhQbuOTrIpi7KhyjZUrtMoXr2cjRYgoyjX3DOCKYqtDG4PgLahGQAg7zhtnAnqCm
8MM1e5B7Pa9zOYRMVZN3GcKmBgvqTTm0lo1kZRCB2b30r0wS1EMXBSsHB2hK4Mlh
eByDq4MBVDGLMFjXMCY7AGghrmAFa4TrnNmIbJenOWg8Y3Ze0qBv1+wI90HQ7Vcd
gGN5pG4HastsKpJTMRzpJG57wsq7BsuqX6LJ6WcbmlJfMBPxfpJAyweuy7IUevWt
eSxkEWFUxceJb8uKppi5uZhYVwEIg+gNaS7kyhpvD2+BEBVDyq5DKafyFrehrRZZ
N1mzcyb/MdbqfFfTJR3zfFuXaYQuVdGFh1ZVUtVqan6m7/dBBAgwgswZPZtDurN+
0TRriCaRNEUVe+wX3K8VSkxKveZoQCIvW74FrU7C5W5OlA9L7Sw4tFKlojn68F1a
b7qfwyu0k1umhLF90nDGufZ+ucx/ap4kLnur9H2M7QyKWWkKg+hK83jitGPrh22M
eHf3HwIm7gtEeiwce8RZTWxsfCofVIOqAOO0VZL4gaLWibylnfv3giHvv0FD6MfK
u1L8xVx5QBMllMMBUNrb07wo3+5HaZVlncabFdzjldhJFAT4r+tlPnjO5SOisoQQ
T2KvN/NZ3eMLY8SQb+aNV4zsAZRbOL/tudVRQ4iBWXA63EMN7d1jSbLHaXgsr3+y
IBQHAwKCcMRCSXSh1TIcdXdqlAlHvP/w8v7zczF2GkTJOGzJQE2PktcXuu3J4/v3
oh9nWxomcNpxAQg6C4eLHGqxQuAKf5tRAB24baE1gq0zZYWvjBWVMGl43YLUkRV8
8tTEgVebq7sAxTtdxeU2PgJoPWKMqaUI4u+16da9CtOReF9IFsREwOlmoAEirHP+
iIpkaUOpUUxkHAqABmKR2+ESGuI7Gwj16Uu4e2wWBw3xm74injeFk5I4lP3JRRCN
IZuxn0lQNpowtJe3PYAEaGtO/fF0YdhGlWdULz/AI44qMXuv4pt70Ma+f6R3sKgS
f2VaTJ+Wxs8au2JmkKHrDSuNqUb0mzDif3ErYc4j0NgBv6H81WrzsygANIreUR6z
z1xOzrO+skleZt6Kodpak5J8InoZXFryOP/o/JdTlJParQ3mRmJR3OVJ+xoUYSVy
EOGASzIoAP0gIfSFK2qKOosr/d7QeuEupkvS4dR45tMNNr9kiFgBozzrU8++Ma7M
IJaCUxsAwVg6+KR0y6nmnJLG+HdjzWkjEZuFDn3/NErWBLy5fD3MoqDnvJSdlwG/
VHpyIL1wkW+oJHZTn746n5NfmNJ7c7Px6Yh4stUMc3YAoV3t+Rns6fYr9fbDFTQU
sG+8liDALbsDzA8TPrREB8/fbODkCRL3Zoa5Z856r6JlC+CtdvbhU6UyiiNC2ZfJ
AFKbd8WASA3W5aNSqXdM4ANeJzVHoWnQKa2Wnr4cafAwrkirhGI9pl4knM7xF0tH
iDrORvWCBWme3JWwqsyvTVZ/+esjtNKohaY4R4I0tVQQVEWFX9itARvm1KJafAXO
wlkG03oYTPjsWeaKtiU/NfkZsaZD3TU/eOpcJHnY4LtWRBtWJFeiaspPRtlNOkWK
5A/C9Mz6z06rDccA96sl+bvc4c9T4qcgTEK0LE1oqkoHSqcPvCWp/5r7rXbx6igg
rgkfnSLUggFTPEX0esntanOrp323nHd5kTbt1VjuHtwRbY3phKo1uNQpF8CkpsTQ
Z/rLRy/En55rcCmSBNBrS2nGAbV2kBLrXLLqyJeXVhMW/GnDr/siKwVLn0vF0ZVE
ZonaA6mNkSaX5rHxrNmw/3ar3rt9f9VQlEAgqaaBqpyg64Cib4m1RBvFTnkCPo5m
mtbXJ7QiKQeW2eGXZFlQyicmrXDbOoeiw5rcr3LUH2lwn1yEpq2JQdkcmrSJU9U3
HtQfI1Sa99l9ENf/XA9A0Azq1cCo5Fhzx5ASnVOdqiwjdBfUJs9mDPWRtet1Q2OX
SK5CdKLxJkT0LI7uwpHhofX9wJrPzB3IkM8SqDIy7DfbNHbPXSSOPCYpZlCePY0+
NGLMvERJveVocRi0cistGBvILE3fKdIngAch9VFwmNlS+Ttm+yPrfnC50UBP+bQY
inTT7S8cOi4Y3A9otUamthZQqI/B9KFCpoF5auTahVELTi0MXgw2JNi4qrImmSRV
/HsWIIJLGXh5aNIdK+bh8rx88LFVXlz52vLs/kRyV8Vk24Gp5Oom2F8tjvh5qgDH
M2N64l6Fqq6jNQH1vMtwayDUZfuZrDKSJgsZS/D1/DE5i4MkUztsFZ5FydjBDo/R
3dhEYznAcTQq3i45mxDuiv71ZOQTtHxWF8KrO+0GZTHxzIX/kWtb3ACNHpG57Wi1
SGndXNKvVQ6vwKyKCUe5Q7NmUuHVrske2JiRwoXtSzhRZFudp2EPjgjnsdzokj77
hU2UjOB+j2e+RUy3ZNQn2IlJKi2uQh4JzzY5ZLeIRuQ04yL6eSfwMDcQHFHj9EpS
Z59ix1kY0lVAWW1RZkDx+QeAAt0KrRrtwSx0p5XjoTwpPlw818qxxg07oaReJ+CE
ruNofIaWsh5ViFPFROapAeZrFzLlIHnNNYatJHeq0HFEy1f2yMoxh1ZBHkCUmN0H
bhnW0JoZJuT3gnu4WdTQRK1CHnBsYZ1zGRXS0p6jVaikNJQHGW4AaoVMffl9dnkz
hf3JHe8VOyaHC+MQJBJrq73NGqbtw4Maxg4wxW64hk+oHFNLD5y7pCYieMG2qt6+
zluBLnHFU+Xx6cI6pgGbSqBsdd1EA9vNvhYI7R4AxDn46uoShxeYmAoJ4dsQ3zi0
CamJ2/z2vjAYD5QXum9nBSNADtHdxg0Bc8HOHWBHGNldoKYUBqvx7Fjtlsj0C9Db
UoeeQualJ9Nkk++BU+FYDZIgPF0j/5E3koZNmhCaAu2WY9glmklnHmqXnEBvJEg1
lXodGjbEh3W68gdiAAzAxL42sH0KKZ9LB0Wj+Cx/X21TIL1lCHnr6AtT8Da//3gP
O1xHzcuQnVyTg6nMvG1f4rQKiGJEroLABonC267G5IaaJIJXujQnTYw45p71sxMx
jiLgHFpbVP9XIiHtSqXutzFzgnBkndt0xUsJjo9GXehq7bBdVs0nJXEQLKpZJ8b3
3ObKIzMRfHA+dAk5YhOGTHW2I1obhFwgfzU2lhnpRAJcHH3CebBptJYmdd0Wlz7R
gof6KhnvvxFuVt7zXOCISYCTeMpqUliOFRB86I4o52MyBy1d+8J4duMw2hKIJy01
NKjiRvR8UHKSjbngCnRhItcYrDpGctRhpBLl5QzGGljrHfV6g5UW8WrAfGypfK7p
rTGhSmkpuLrJsgS6jIzBYSgHnvBb3cNzdOajsKsdLpvJH5Faw+FlkHifCaL9zKUC
nbClvsS6hMB2bY3msYrhupr96E1ZRKthvu2HOxPOLYHGDNGoYuGB9Kk8SAsVRclx
yjqa5o2hvqWJmqo4J0+UHSharvSsv6HvvHvFSvTxce2JpefMGpEgXaNT0EENOZ4E
1VxUOoTJe8iJr62DKN2iDjdcES1bQOA/vMlmo6y/fscw3w4RoShvBPuck3WMHM0D
zEGbJWTdjadqgu3S/1AlsBb2TEQgsABDe09ZguByZP1JlsdaLqtZLpFT2CjArwX2
GMXq5RJ4YZUJqQ6axarugYjO5qNfLnrcVoMUpXNsV3QWZGlcNDaTu8024liS34Nj
KtesVb33bYOvpZUg8pREqP09A64ZhchCFjFFqmD8utptpAw6PGaNM89irHujDb2a
gKox/2r8+0pYr0obZT0RuJqQOYtjOxX+GWHimbC9oCLi7AtVM6ZBe1WQLnS/dUXF
b/y5pedgfllnA8PW5ukr4hnddZfG99h8Zb3R3+2edj5jEEBtcTz+CvKM75qqJnzr
/HDnrcjWwnyQpEk1h4rnRGORrE5/fhsyZduARWsnel50GQwwpnYZED/4LsSkc6A3
CJZPVz207VW/yPlWGVkt7DAAvf9rhu1D3fFgjrYHVZiKIX3gookZUqVzx14PtLXY
BPEZc1WPceFXePHY5x1XRnOdBzAvyrGLujiT5Nj0vqA9fpr/KovX9E/FmBBpQ9n4
PFEfsQwgzZFft+NTC4mnvdTUk+5eiaNq+rzDTgLIwowpm0C3hbuXd8ZmeK7z1ob7
qFWtvc6GSzLBzQDdMLIR1etFBNYvlFafEe1BzKcIH4KLbzhsZCqDl0V/bINyP2k6
viNnftxZHxNwWKEKL3MHzHQhjiv24Axa4uOnmhox3sAq4w5woRRh6ZWGrfPBxGjd
IpLUhEjCmtfCgHjUolFKuNQ8ja3FFS3N24yqta+LOOto4E6uOPYDindbSOZRgEGn
S8xHXSNlQO0/Aze9vHcQtCXqhcH/UoYP5baVT9k6iFoRsIVnE9HHGfHN03l0cXNJ
n2bNoKvD9VhGEFdbVQIGntVo7SeyRrQhM/9GJ56mJaVnPAH7uz/7d9IfMnEV7Jml
9QbLxsn/SSz+wumQsFBzHdcQvnAWMC9G7iAZP8/EIHZE9+6FYLRH7vfPbGRJaDeP
GXkWXiozg4EvDXjEMlH+4UE4E5jt9GRzr6a6k6DeYg6UIW5yDCvDhuVg7r13olt7
YS9yzUdv5gRMa8C3wNRtdiYVDc44TM7GztlIUq/R8/lwiV7Ghg7b7fGTwgjMiowL
P72jfUltmKZw7UDqB4yrQB7RSP5HwcUR3RgIs3zd08R91B9aL5i2q0YL4rYlnkOY
l3GzhkQV9FIjB/13PvHFHGWc4CK746Kn4jYhqICSTiN0wE9tz3aFKJNnk7F6Nkhl
Di2zQhMi5OcnMuamtcxMyFe3XBp30apw1s1aI3sG3Ds5Txw+gOKb32ikaUGMrtdz
C8rNY4ej4OjKxdlr6dSgvogaEHFM2fV0eQQZzOYpV4glMl5gxbWZM2XoYV3fITaE
XI+VRFhe2CFZITDzdB7mlWZYJp6zWXTghvC1vmGCT5hL4NQYdugF3e1Jrcy5tDWf
52Xf62rvxuSjEIPHddAECEEdafx8bYHQdTs66DpphPbLZnNblZ3oIiPDPhwScKsE
cem5+wUMNRrMz05qy/bKysmW6tFgVUqfAn+4Emu3mIw912zRBrX2xcxMdo8Z8Oty
S9mnQD2yeLR2F4k+nM/wW0ZO9aZBDN8Yv7BVspnviV4d9/YSox9GGwRpQIAQVdCK
3twPozvHTPtNgemA1FzXYx6//dPoxHcPNsb+/+ZBbloIz3veXYXXD4gVjYCIp8hr
Zx/LwV+1wZ96LJfXPbGvyfSjwODDd3lnqE89SKQBXsBtikGOTBRLRxDYqgfCkXAw
FKihlziPAEMybfKj8ZNJpmK577YnMosOjXLQgbvO4SqXxNYyXEspidT/93g1v6lv
snBOqrsF8W0k4C5z8bIqaH/GCZ5YVlyIjPRggY267lPDQ0gWISeQ5bFSENLXrmvD
gU0NLVajKYAOMbM8NAmevH1IRMbUaBrDIQz5We2Cc9TfBhOL/K83c8XOLb12Y+7w
Afi7M3CkuvApW6VpMYCodrrEtFsME5h4qkgKsdFr4w/qhQpVOFLk1v0Gz0c9BVS2
pF4cWoANrDrfrR6Zge50+mBVLBGZgfQVTokQLysCMDW9QjfIr+ywMtbIFItSJ/8Y
rWJWmRrWQUWk07jkeeoSPD/lgsVb2AxWrDnJcSpp538j4yg8dmC8jZf9JYjRALvG
UaNYQPw2FVnC1g29qazlrgq9x3mO9aNdHgKjnBDzKNphtuu/3kqtSDRWJlbykt/m
0f0OIC5N7xSMvU+8xs//Ijyh5wTpdigmW5I0QNjgc1dCsNdJg076nP5gkBtgk82l
9uJ+wCWVjSPF6dYt27oZgXuTMTyRXX+6Skv8/BUgx1IGuqOQaSBRPZzS9V7BQ7+z
MV0yBlJkgC8if3PTHzqx8PZ2hG5p28wlyKm76Tv23KDUYzUZ/8T3jooP10gTP9Nv
x9Cx75cYWEN/KpbDfYXO5+Vz0NUeYoxYGvHJh1/0lABnqojyeV34rjT9+ipmbiH0
oa1gp1E2RQo7OlNy7dcAC7fQGK1lLBvYA0MlmVZ03vRdP0cldogiUV6pd3xcNPiH
spzyrFslUVu7yvx3dzvQE6BWk58y0i3XupMLdURHbweG5xhrINEGogmJVFKQ4mxg
aXUTZYn1FYpIjeu6qznngXwGFqhK6gxu5o9yF3zfNd7KaVMSDJhlpp3o1LUMpESl
mQCqlDV9tthWbhRE5hzmGPH+TBXfeW26mWkLT53h1o7UZSGBnNfRyL8LPzqXkN3g
iZDZQCXOS5arsBf/3HHAUZICwH0Sqnw53z72eICVbaIMohQ7myLCOOvNMY9xQHBf
eSq4YKjwY9s74u91z6Wp1I6cpqCKzB96Rml/Tdj13iYXwIa7+wJeytWiGM6pWyat
wgZC/CJuT7AOSgCfarAOlXVoG7cGUTJR++eJDeHQ1JkcvWhumEjAmA06CkUgnxph
JsyPQphRYsIWGZQitL0SmrOcCu7JWd13NJRk4cwrth8w8Sp4VQUpXoDr133cLo8M
W0DdaAEvOzbIgGyPjJ/qslAjLypwShbC8b6JLbVqdAFVjZ050ahM4nK8Ia3Px3t5
W9rrhu2njd1UHgS0t/Hea4enDYDFL6SL1k28E+V9u9cNVoQTjOq9HCs8dDtFq5Sh
qNYLLh8wZMEQq7TGPfTRbKj0fvGPte66Hf5bJVCFkkg6av5q5nfZFQTRWLy79gF/
yToHOWWF2O2RzahATIbDB5AAfmb7t5gOoUhzfiAjO6vvR9EcqP2+VgmWQyPcqCEa
Zfvp36xrhHyVmgi59QidcpsIk/IrV9LYs5N7gZ5UcaSvIO3tpKgjmMZr+Qwl2N/S
cbytsKdRFi+Kwy2/bd/wpmJMz1f2RA7QRYpU3dO7edL2tVFTV2spEjYvb3E2l5i9
RxHRRySVOHcBlLJcKvKvpjsQrnrUhEyaP1mcn7lbRf2F1BeGyWOgQv555EnW/Ogd
o0HmIOvhaqfsw7JtFbioC18qu2PVxbvEQgdg4f5n3mg9xayAQ/YfJEHMJ2cy7mGx
TZGbbmmzsM8B3iisaK8qi80efvGHwddmL6RLPuZ/BDNU90fpc05pU29M6OIaLYjr
iSvZbiSYXMbR4wET4N7s7jW4YGyR/Z3ZHbcw6zzpttCNsT5HJbPfja5xmDQEjGVZ
NsTKP7zz75Bv0zU+7gbAKdlaT6DKGLFx3ak7XPlsqfHIfKqVJrdwuhAYBv/zRy/r
Ozlheb5lWvW+GJEGBCxWkmR8s9eQHvsDKe9o9Nq362HmWgHnmNv/RMPSQKCHZ0SU
F8XGtzzr/BqlEhfjbj9aYsWHdHhfaU5sxhsQS/B5BZnuAUqsgpXRkCrSKbSf6pBe
vCesPr7za8jia7DKFeCv7+l386tOA+yGxcuVI16FyQfsrjxFtOcFTZ/jNKQSqD+2
sNgoVbpl0Lww7h+e42Ef/TJaBcKPw47KSMdC0rxQ4gHlEop8/0TBY46OYAlDkz39
xPH+181FKThioj7miRgPzfZlw+JmqAgD9c0VBxxc6nu+TBVDvrU4S0TScmn2hiUu
NPzG8O7Z0ZcUA4n98XF9etYuxXeVIUasf7zXGMJappRiW+t2HCWIu1s0DIxw/l3X
2GBJvInuH3LzGGfLOZf8TOmnzVAZtwEc5bVMax0rLncGoTbMQNktoCA0+7/WmEz1
fBieTc94Y8IYKt38kbUmUQ7+xVGcMID7KP+tgY96RvSAxOiwYWTMY2gpf6Smy7Fn
JK30zUEI76XHTOjFrIT0FRafvh7pz1PdGr0FTfPsXaEwzCHGP/vcPbRU2XU1+1CO
bKYOUSq9tI7nN5NspqPJHnrfLFDZnZXT3f+a4nVmUfjQ+7Ze80PH5SGbeHZ9myg0
DlNAkjItkTS42kN3jZvkAY1afKm/oryPPFaYCxnAchU9SxdJ2qczXN11+qqNxjeR
89WhgHlrpbzfDPvl5OlbNJAl/iYFtozUwMwU0WTgj3+Wfc6ZgFzc3BslNWOd8kHQ
r5Q+vPdE05fpJS27oLdQAqz19NTw8E3oeherYvYEtIq3/M8gKpiwZ9/tYZ76Z/Zm
QMmIoM0eITF3WnFx4q8Ipzek/1lGr2MBmUnKO+dJgArATMKAI5YYsG5nAta1rOJp
B5krdpJb3V7pQJYjPkONjyTn0uetLm4DuvGOvsIA4Qri/6/sAd/H4pJ6wboTwQ6O
lkj2R1Yx0BP4j9hWWjwOrNFM3uaMJr8RQleisGu0BN2q6leWlVTdQL0D22Nw6jqU
+snR/y94XUjQKeD8pUJpCoozL54C61Iaa4JtkbpMAyut5oH2CCduKKbAcSDWvFIt
N/0+DyqZJYd36vuUWk3tBUXeQxX42QaxRG6eWYiKEHHddK31cIYO5Es69iG29Tuj
p87X7/KvZvp0LbnY5YQpE1VAdKbjvr1xgjiKDcXXmTEYi1gR8fttX/kVr7N+equp
BpSGu0DlNg9eJTnjQH6png7mCGD72PRRzSySUTFtmWYjQh6mx8UnvzrvDkPIzwYQ
or2V/5Y2Ye8St4sqKA7DE/4626RC4Nq5nJe7z++tuyteN0KZBhQj4EpVT6hM1zZc
vnPdtLbI7/oNvKucQiH7P3PVRIBLEPglczzc/HHgYeJV5ThOlWzv7ROjRg1BdUVv
qOdCeuVas5uxfLoKJQDsO9ANr/wn5zJffqMkeX9rWkb5LC1oFEIkIy5iQ11YnKPC
3Jc80nKfkxduU0uUUmgxkuJhdgAeeSVILz6lJKCXvGL33qBRwZKdi1LUHQabQgZY
i6G4ajpieq/Yj4SdQgtdzlERkjqKRZ564dlBSXoY1L7gBf/caJX0dk/KSL30vGfS
mK1hq4xYypOsuuWxNZlXQVzvQJ/sPn22h4gmNOiD3amIxZmVH2vp7k1+ACcV+2V/
rU4MHQNAXOV43afrpNbtMtHH2bbdrTPUa1VCftsSMjf6jpGq6ZsFR9HF2Z+tE7WR
0DjHF4r9WlKw8lXuwTY9cY4aQ7Y13Gnn36POmAykSi1P+c8hhmcSoJhrkLUbfUd0
BHKI4v5UnfM8duNx5u1Z/KqtrEvx4YGIDI7nqNYBwxBd8Yf/F1L3R66xfjTlRsu0
Xn+d+C6bk3W97vWbQOVtD+o5E/DbT8EDMj9esIJrwvZKHb5Lilp4QgyGc7XzBsUa
wFv7vlmk1Pr2R3Nd9lDOShHh3jEubheeYHl6mXlea/CbEN9mSFdvZc/I4TbOnqFK
7siFaiV/LPNzyVVQ0Q0RAGtP6Au3Ot7c6F5MuCG3DU3rvn84qrT4YkVxDiJlripj
YxOgy3LtXz7nPLYrhckQkMfLbHUG1LjmIhO+Z7RRYkGf/et86PUk7Mk3wdU0bU3W
aTccYm0otqUXW/uDnTV423P55uuUqQXuMJDLmAntYqz+FGnQmUEfPWx1BUX0xWeu
CUt4qVjqQSDoifljzz54NJwuTsUtlIKd7NL7AfAMzKomnuUR8nkkDO7jyezM3y7h
6SGOEsONkt6YEJ8/a6QYNiKd21mQRI+fuZ9VJEe0mKqt5cK2M8vXA0XYqt1+sGiq
vrYJfJQsqY+CNnUKGGOm6YCnsvUpeRRJGv6KzL6gFpB5G9J4YeM/BydWSV8fD1JA
gqsYef5WVAZ2o9/rKhc0tHWnTX+XA4AiWRkLtDsoAP91wCjqBx2rsq+j4dn+O8OP
3LI58sPWccjvYckIDlWiwr8gLmxbsv3RKuWhYiaBo0M9AaP/5dSoHyjYO85tRQbf
mc0u977VcxwnXMJ0qQ/ZqHb0DIUlXXfAcr123pEMss3+XCfxBay3ESK2MWO29Xy2
6sLRdj6goqrOSjXInI1ZDo8tL8zy2CnGy1pUn7DaZyJ0vngUwOSFAjTTr+X8cnk+
VF/YJr915jFOfM4FeAtKsJl2CegNrmGRb3G/YjgzIGcMLvS1cuGoxVpE1paeTivl
baMnIt+/ilrK4crSYHHCnkEHeQeQGsui6gyVyUiZOqBc1g+8gsWF91DwNmg00Fv5
bB0PxCoae3iNmSKgjYJv2cIKMX0twKPPJiWlMXjrYxK/pfsxokSbzgI/WQA0B7GP
4EfRJYyB/EEaD4A/adbbVJUke3KmlOZ4fq0i8nmO3On+D15iIuHatNHDc8CVeYo0
v9pfwGVhU9VDT0wGylPSiWSe4eWQRe2/awBtJnER5jCiNLbYrIDr+cty+0F3rvgR
ZdIRL95xGWMWk9lYGBYYA1In6noD1H/8SfOmFlwPyyp15Ue/+scyDwEkh0WpHMVW
z4j9AsPSQmj8dPu4uxkNULFSJOyDm4hGXqkwWU1HZKDy9m8A0IJEHbEo6YMS8erO
SgLZ5BvOJnauUXUMjycuekyTZSsJKF7t1AwqMtjk1bJUHqL6pl2rACQiiPc/YOAH
OYpkwIsJPOnHQvor7W1WyssJX6P3x1YtJKdxnozrbz9OC3l0eMan6dN3u/YSbpNt
+3sUnY0xGKd7OOg2WP7czUap7I6TxPN3AuOPhqFX+KWumfQKwSUwb8YXB03Yh70l
ddh/9Z6YtcyCggXMie0Hr1cFv2cZ5JUxAUnqD6u05ObQ43WhOPbKfU0Y7lNr4zId
i6i4d6dWuuzZd0vDYv3wcRD1qGs+yCGe86op6Bbm0RnmP9pdfQKYpHp8fvwq/Lkp
p7v6b9N/osktUawMOVHlrosLMn7x4PKSkIVJyCtrefNAMT9h/Y2DdG/aHvIvo3TJ
wMoTHEwkq4ROTuojOI7zioMG+oEs0vssV4HobepO8g0YKlWQIk1swzEEyDAzmrz2
g5it102wiQto6zj5GQSgMomTpjzvG60wNYEnvtSONbJmeOF2DVgENrVFFAujZXFD
6MB32KQY6DA8qlTKlp8y2xgwuLwRujqmlxYbWHnyVwQ/eiOoL0CSusCIt70/nh6L
zaQlGS4OHMDY84w0QUW3v12DR7KQ0AJAsVCyCEkvoevlctiQ5HWbVhszEjT51RM+
W8c/EEiyWUgg0GrF/Srz9lNSRUAKpNr3mZOz8T5FkQRFMST9DHpfiuCy1SNyXKS8
7Cd6xa4IpiiFmM/f9SpW+OfBsanmvz5PzrnrnAPwziFOIXSPY2NOvWDMWyoFrgl1
LL2KiH+MChV4QcNAZvtp7Q3dDYtPe7FjU3zgtsiatcfspqgU+oiBDGIHnOxixp7w
FnHtyHvqZPKiAczSBr+Coy69uW4B3gzTOf0Og36BPhg3kqqk23hjUnkI0SYWg3rp
Td6qr1hRE7Mh87Y5s4kFLvPRgp7ul0+2ZRn3eaSUVF3ZUcpjK91Chj3hBHge97Uh
6IE6QvxxL23aU9tU83GbxNvSMrn5saP9nDFXsASTNvacIEWjLKnBAwY0X19zFW7D
SaCRQ4LAEwVhF3749Z70VxFWhZzcdnYxUZcC4Kax8sQ0W4DFGjVfrMkvVjv3Z4VX
YH0kfYvy4PPBZ+C5Yj0nXYsNR3E+nr3TWFQfjb1KHvvNraXxv9PDkei7+E0iAQuq
0LoEOBe9cphCB2lyxm+AoIlEw7WNSJzyqHopAWhnuGg/x8BwSfJfpC9cGtTH9vxn
OrVXwM4DTL29L/8as/KkUGqipD05MppkHrq6whRHoskJfaCm0wg0fX08tf2lXLTU
ZwPKQ9dpkks0Y9P3e0xM5Tdw5YiqbjIqIPjsdcMDpXd9YdcTCa26h6p/TL4xz1R2
qHs5Lbv8Nr9JBsANFecMDeYcyqwphSUQIIyOlW6yLcjx0JsARkSgwKClyvvFnE6v
AdgaRaKRMfoS3ASmNaZ8GwOITj+N2yhsyiP1r6Ff46SCqaYP6SGSRNKPvRwZrdnJ
WTbpmQPooy+mVyTinXYaRn1zouB3IvzehG19d8EHbWmO+MTLVzvsE1Kaih2NOes8
VPusK6lhGmvJ1xaT/r4wAzqxQNqd3FMSkQCCkXX+a/OUUaxkmL0i6DzBo1E2rjRG
VraQNLu+ruoMyUv91eKD/g8w18NDEqzCBF0e1tFUAUfGH/cUZkyji+abxyPLDZy6
jyBVPgtXCLrXQsNG746SuxNGwFmPzX7Sw1Jukb2DRCx+JXoXVhdZ5hJ2o0MqIa0h
JrtY7FwVivK286rFzZCgKznbWLqVVXHowgc03rWeRAdL3vT2TmnT2B4deqkt3/pG
ML6cJFTmgJMciPpsDG1/mEpM6+M/BCbuAxPR/ZxzLIQvsQe8dimBq8CGdjCn9L9I
hIkvFZ1rWkvhgm/0+zRtYr8fztsYroWFHO/15mZTotnYxLYbTV31c0nsZuQbCKUA
6SHB3RSy5Y4j9q62011vj2ifaryhuZ89jAhL4jF367pw9W5u7CZ0ASEeJTe0PJ/5
5KqTgRaMRbmdqenMYSzGaudIBstNtfDEewVptL8K0lZNyXpY7oKSqRKOYrGQHcWL
NFOcqtRESKjj5HY0UFCKaJIXUN8/C6hC68uimwnslHl5eAaxKzSCuioLAnXkZToS
q4tO7/0C4AI3oa+Wvkr/q9AfIiHb/kH4GVQD47YZlQ+A+qbzULD5k7In2UIPeX2T
jyTYUthAZrhXo0ZSh+EHUrUpO3xEgRpBRSYDROwumjredZviid1PHYyMYfVIiFhr
3qSNQrkxLunDVJzZe1WBKK2CBIh+R65P9h3qYp97yEevPbd0dnyYMBM+dzJDMPiO
2VLOlVFajprOmZFQXFKBHP5JLQDOz/JfHnlBjAoGWj08nzFU5SJDjdH11zG7Tu90
j6aezS297aTDRWLzfDnPL7Af/Dx7JyaXmKxwzalLKuGY9pa3oSofOz2qZ5xp9OZG
7zitCwx7B1BPq4fh5BclRyO1qt7aYmUktz2fO+ikIy8yXiX9Qu3RdPd9lqz3Tirn
dZWM+8ALWYtDlssrPf05nFBuEjvTR1V2JyqcF4QWlbZsJVWvE/odGpUErFl/rL9+
Ar4lFc8G4LWdmDuzU6v6piqXWehroCzUv1J6y524hXmhFmPtUDxjuiwO0T5mx72m
MqFiB9AtDD51lbgd9YC0FuqPGhCmHFD4TfIlO/aM9FdWP1p5S55MuBzQdSjIyCcG
EJoPNwurlSA/mws+1QNIX6CN+4NN++X4SnOG7d+rBOarFyf4yj5rSGMx6ooujStP
EZ1W553zVOEa5ijV8yVxceIhqMctJCp+KrZZWdpvMN7SouxQSLyRaXKyAFDURJxh
kYDAs2h7J0HkcEOfBYytdTYCPj1tfdv6yvXR1WnJu+rRsV4RXLNgoCiBgoKA8cfq
SRmfMpAwxUmkyrNWxWEQqB5gMaak4leoB6VW3FQyNgVR49M6dT6/+qI2KlQX13sd
SRMChtkAfZoyKjpi/Ho4iY9H7Rk3Mk9Nof6SUFtI3uWk5Kj9Rv6f6lj8tJAWyXMU
JDOyij2QwpYMrQ+d2wOF+ts2jA18jXIe30IIV/ZnCNYLGl87yl4jVUQ3UitQaj3w
nvByqN23l0uCVXUJFGy456+7C8bMEdPUFt1uF+PH+7riiXX4cI5hqZd3UG+ZFfHm
KVBHWEqzhs3aSlAw1oQqFzfWqjknII/UBv6MGC6fa0goWv5v1sKqshFPhnszEh8G
vXa2boxBiwE/kdzzggnzuemPFRY7Rguf8QGsN3pRmJqBh6/90UP0Vf1mw4mgnmS2
dIzUqdfvySs1RVzTlb/1MRZCVpdVnDmFFtCp2YxwkDSf6Dq7A3mp+VImCaEsAHWl
i0+E0gJ+u17u+Ldvje8M4Ync+L8XnSyvjX+lNkuCyyL6e0Dog/QF2pWiNuGhStT7
cCd34UaQ7kdXJkm6F2piH9e6bm7nyuhCQnmUyYsXEGmhXERPSRET6pUK216Bvhk9
r7/Sle3sviIeL1LwkuSC58P/n7a9XeX7pHmNFvpSbrQt3XXMfEOa63v4FpaZRJwC
4YnyiiRbFG9X+bP7aFtG8Vnb4PpNKVLty2lGk+TL+BFx2oEWb5YZBCJjE1w8dvj/
UJDgcxRCClpXakbeivxfkl858vArwX2BMoAyVd8xZX3m8VXs3yvjeZr5AUsetqfb
xlrZIj1WxRK1U0qLAiIDwLOgvLcu16TF+nni9yuKMdcoQ3DQprXfmt2F3Ak5OUOY
JHclqCA6vadMvIKRmWi3uZATpApQZj+j0WmIP/6XhowizgFsJbnAC6cEk71c/h9b
k8bkdT0jZ/SRiLK9zKhzZLpE5ebyTfStfb+cJYZlP9nHFKPfXl/A559cYF8Nrxk6
+CoIKOTm78PiqbJ9spVWgkbNyh6XgSINmZzg95pLczG+Hplz8RCc077T8chctQT0
z8eJo7fiRbKkJxjwAHWoa+GMg1YDntdagobv43DLh59Kl2pE5zowlFTRX0Rfucke
C9OI7pq294bXcKNWpARB+9QZSuzYkZTfjw8JKzNfi+DdDPIt39zY1WEs4Be/HIqu
rdjc5ImUqdLu2HlkNoV2ZhfZ1gWCJ9V0qGsBHkhNn4ICHxjoWvucgn8if2paRo7F
XGDYOSYAp7nrvh6RZPeBwOQxD92Q0I0DO+2NLEvG4wxGHYOmHjPxUKLwkZchcD03
G3qldZadFEPhVCPytUEbT5dlVNBNYH/KBXhAUqtgkaRE/IvbTMlwBFPTHsV/UcvZ
nAOLZT/vbqJzoOP2ABrzMIg8xpGat/tHSvY109F1RXBDLqRUHnMoi0FfljsWjVpe
LOZEY0OazyXwBwo5fG6FvkvRedySGC9kndqa5URjjzOgg/qP5eOjqYktoVk0m0kR
DIx1cbjXW//CHwyLNVokjrtJEzM4651pZnXWVcFcmwGpFKWR8yRdQC9AMISu3+Ar
qc4uzabJnunU3Nn1LVkXkdi6YdOvjZUWeo1CY54yxc4K0kYyowd0tggfyWqiV0/y
DO4mo8cmyQbaXSVMdrj6obeWzdv9bNC2SN7RqTBYb6dy1eOC9hTXUhjlaVMTvgYh
o0aT0p/P9O2neskU9ZBnjrAfJk5cwMhwKNC7D6Ez0zzcJM+CD9Km5AhbsuHrYgJq
cqyQfdf2n3A5cqunos2lHu+rZJyrgMGUUSaYt4bnsQfkjxZTPP/p+sFso8TLzt3v
uyVx68n436ZFISOPEj7r+EPLsphjDMGW8DFc2IDnednVGeERtQaHVLjigGw12r85
VZhihgIpHbuKO+JuMPUhtwI7IJl/iFaQ1uwyvC3QsC2CBL2SAh7ZDibl6yadGEMQ
oS3tUnjEKXR1ZQfpI/1RHMOto6x6NBN1ui17ktqv0XYWViSfAmOdb8Z7geG1awsZ
G4gFs/xz7I5j9CkdRSRakV9CqAY5KW88KsmUnc+qCuB7gPnLjzZOE5VKaUSm1vc4
xBEFxbH/scfA+s/iUb0iD4pVJoSXc+95TCatBtjZStzngCFs4l+hpY/H4yA7F4Jo
UaW6jJzV25A2hEOw3kPFv2q88G7Z1aH4B0yZgztZfg5QYPflEtagSGVLDTecCKJc
8wFudCFInEoBhxT9tBW9iwlMbrjbO4mLAqN9Kuos3CqaV14N+jiWE1BPzQPMhKpm
2nzQ31Ts4iORhI98xHmr3RsgGYNWh6caHFvIZxUlarW1oHmSEOnxIOA4RKw8Ov58
ahu9HzY4rVx1VkcR1cmpXs90UggKYnLRLK+Wb6IZpy/A5d5swPHcN5p+WYzDjcHp
Myr6vkLfT5ODfuGYiiJmoiMCKZGTMI8y2+QREGe1aoSp93fHuR+4VpEN2rcggeS2
mVp9Dzmi7lUzF1uoKnyzrnmBUtnN2iga0jyh2IiMl7NgRiPDcTKsIhnqD3vuK4vs
reiYjmJB5vS0MgzsIRabDk20Odt3bagW8La/C8vAlolRzPcGEB2PaiQGZLNVqoXe
2qtSY2l7ZP9EBFbU/8YxHnP7dcWM2Q4P03LpmJHHHAkV2a6qHDOG5NoN9/ZPHfOc
NIoeBthuUUe9P+6IBDbdEeiUZjfyHRA2K4n/OZ47XK1ckSSg2FANjZQXQ/7foEXC
MqRNjjO/+/1byiSJ1WxaVfjq5SU9k372qGPW7VFFKsTJHJ8RLTRrEuNgqbRfTMab
3Me8vpAgfc9QlZo26DXIx1I0zIVP/OyNvraQgpES1ECoaBWwUpGJVfXX58t3VjGZ
MvGuV2VWwpLqOsM0tzM5GfdW0bKjSOKlwuJxGlbXeliZ1CJ7SVgTeA50d6mbp1g/
DgupTL3jVP5Dt6C3m3WVGbZk8cgb/oFcvmfaDXYf97hCstRUzAkyB1R01ToeFsVc
wQk0GMTeEP3dBQLqmQLQFl6rq6O6UAzgwIIJdJJ1ykYA1+F9cktSSIP3r6Xz7Irq
b+sGlkuu7rH4SdV76Dqpzf4O8iKoWQVBUCQAKSC/fVER7uFpNGDvdTFyHGRuopgI
JEI1530ZfAS45ZR08A7S6ivoHVJCKUBc423LcDVqpsgi0kHCQ1iS1ShQgGPe60I+
mUJUPkKFi2DqOvMT0gw73JM45/iAuCK+oVgzWspKbePE08rDlHZeMkrLrcne6Up/
FKvBHUCl7MxvDxETy993A37LrBHVWn2tX80IXF+WAPa6j2DzubVZvXOLsDb0acvG
Z6dFAogl+sPJwmgl+c1AxEk6bBNM8Xt6PK+OxkldE+fGO+MgWyQcZuL5xT42cpgH
BjLSyeNkEIJGxp7rCKyoXQhinisKf64TKK2gk5KXZGWNop/TpBJl0HSkIY9IR/Uv
EWcvMH8FF+tHN14nFhv7ljAiH+G+MgCebw2RcTu2hv2+QxplI3brWqrMn5Sxj1re
0lvcL7W9S0DyUIc3Z0uCIajoilm04V6cx7oI+vy18kgfGwXzOhMaWfNUYx2WhTjB
JSXfFGW+u3W+5UxdUzIr47n1eCqIf3DjT1iz/RWFxJP7fGhYD6IndZxeOtnSj2LI
1boTauR8t0LN1gOMZXoZVQf58gBO8ZORRoY3Iuu2Ryx2mgNJRWILftbfuz8/54E+
zIdo0N+nzugrWFBvkVl7RJj0KxvWrBDV+lh35ZRdiAmCjix/yvikVa7u6n303QOH
rzzrW2AXX4eyp1ARqi3P3H6ddg1zhusMdOMCHzefahdb0+vRNUScMQrG0WbpK2zj
Mv4X8AhbXv4I8bkmq4o+kPzG8qolluqcwfbmukcmvrAcZTJKvx1tj2RekqLgw5bz
HLjD3fBcPwmcarpUoQwz8bpjsI7WaISX47DsAaEcWj5pB7bY+gUf9r07nnXzVv7B
xWaS/1MM2OO+ezA/5hY7fZDf5HeumO8vcQlVldLVyLt3xdfRP8hR34qcZ+GIF4wY
4yVjQ7mluiMfniJLJYQsuaSPyYArLhWciDzADjR7q54+Ls2I8/GcLv41RrBbpdXP
3wBS8NXHNFmiJq2LICTuRA+gC9m5C7Mx40ymxWytQE+b10Si02Es0Mc9WKIWxp9S
sKx++zy4ZZKhDCucgk5cgSoL7U42jSu7JWWV6HlZSOaj0I0dk9NParND1E+KOPbP
kY2FW0ljJqchu7zvJZG0fRXxJQXJeUA55liBR09zzHg7N7zF1yzfBMVb6d6rWnek
c4Pd6YbypxEwUDpRtK41BW5ihXtUpMkZcHCteWme1q+lkT46SAvq7ElEt0M9heVi
0OJUqY4DN7S6kvQlRGipjOo0EugttM3pmX650RIMQUi66lRwLIC9dRrIwlhhZsLw
tlNHtJ4RZ7W1vIEalqK9UQSz90cWZu6I6iwAAA60Vsr6v32nnzW1NIQqn7ZW0GAi
nkEgwN67KmFCaCt8khhoXyNPj+JiTBGftC0LJNfKBt9L4qNP/sqh184IFf2OBFUW
A4Hb9mrbIcmMGLZQ7PPE/EUrQYh9t/6gwGr2gdO+lnVvqX+qFIuwatWb5HYeI0Zk
LedFI8lZu7sQy+dYBWnY++PtTTEpKgyD50LdKVJc4JZSt0JU8dvxcVCOlv7dLFu5
Sh8aXwi/TCZv+0UyJHOHF8Uer2UDczZtIGPjq21qxGBhZNe20ZcWfwZ9iiFTXfXT
DxVsgy4pQsZIDo4p3aYd1HeTgxVc554wQ95mtGG3XG5KNKU3xFCjT7Q3YHmUb4gg
DUGZn05MTrk4/qQgPmOuwYU3fD7JW3R5S7yhpoj5sjIHCjQkg7pRc/SE/CVxSEks
g201MwuLpVD12DBQcCj5Ooq2f5ACyPJiFhPAhvpXfeWDduA543ojYbepA2vrxr67
v0pR75vFszjbvW7tYCR+HJS0Qxgp3xZMCoLz9flNw3QkSYkeD15PA9i6UnVjwAwm
VXH1vAVt+7dftLjMm1AdH8tdErcgFgi/ukgVT/Zv9lMesbw0IeC8VNdMMsybjMVc
zM7LRzoD8iyJxNjVU7EsWUxuNukBVUZj/C4wocRpsGgXhRq/mHcLsyfroJ67GH5+
8JP9foFSPCGCo3EC2A/YnreZ/3cf717PGn4Iw/nSpKa6qTMO4MnJPOyOEdOlTQky
EZJeRtcpuVKjpUnJNJkMiXzVc/xgTY2FyTigY7r8YuMafQ664vF1bTiRsXfGb5sd
BmoZcoh1JzgUjSe4cjSpyhSLsfu4bcRhXbcbajT3qF2Y94wIjz+L1OC8TUxaNGRJ
K4rXo3itpAUXzAqIOThzoaZ95/3PF0akyVtl0AelEnzjaUZqczMzGCtjgeLiqOXJ
g0C+P+91MmfzAQo0B23UvkZ1TDIBU6P2CMirJ/562HBRJZ6WOYTQlKxjWpBYdfVl
sY3xu+zRUnfvasUIAAEpx8Z6bp4IdZrJ2MLZ/sGKMybXsT/r9JAtU1zUJEPPGb27
O3udCvtshfzrFeR2zcbxZBxxnnQ6Pe5K5FwZEIuuONbhOyyX8uZT+w7ndCuDr8Ke
4GT24KInDt5nxOzcmtTF3WDGnftJt5pgTryML3HVTglkp7pey5liYZHGe+b+PlIK
3haxWoCbEsrtcEi9jJ3igv2sS97CIkXpeBqmkctNCpITVLze5TDZdrIb1ymd+CN+
25uO9VSaWMK6cB2+H5dSN5qqgEzOGr+cP1vqEV3TnNWntZRvfY0YalyyW2lINQo4
CxXGfExMB4897BXFDJGlPJt4V91SH16UzHucANwTvBWBi3vikpqWpp+CgNC9KA6g
9voDE2W48w5frSjb3Am3u23mb3tbPrQ3rMhFqByfZvsECkSE6/2ZK9iN0uGVZJn/
wyDZFH68m+WbGKm4eSZqgGeJjShg5+qA/0cbAX8CNIWYjh/kaw+yiXP6km5EY4Nt
vH2i/C4j4RA0fscufQe+h1LsTGKMnhUMt1CUiKrXoNdgugvPCE6TXiR+xrZSxAFJ
3GZessG8n6hbS/bQZoXrOnCvxXH7L98dfNXxG9TwdpoLYGffp6JsDVzFYd2xAD1w
L5cq8gTrarkn4nczUUQ63jvaYGURfSVdifZIWm0L8O3pRLwmRno+cQmyvPERkcxP
NF4yNQ6TQR1J2O4BxU0Ug8MfvtwfNOf5xUtqM5B5VfnL+qmnnsiW8cwvsIU7JR3b
1m5s48VQ9NR+PzQcfgnYto2KpoVC+MioiiFDnJIidpMOXTtql2yIp7U1Mj1PiwXy
TuaPV8HOoo4f6zBe2tPl5L9xyrl0uJq5WCq0WOJCM8G6bJodB7GxET36Tul04Ik/
F4qiWw9a5XyZdjXrAaNDfDaPiIgeW+muwi6AAUxOH3Xj7m2/BWV11SXfDFGARVM4
e+HB0Rgj8Y0b7whzPkol3URMDEuxLV5N/5315Ew3KoakR6FkUvtp8l5tJfHr1kw9
cO5zm5Bnxgs6TSxGNgtkGGST650Ze4jFe8iNa1DnL88/t+7DaFao4pDblyiW+Quq
ET6CHi5BTrpOunpzDfiLH40rZvq8NNU8tWIlTz/320vh/jHhqRnCtItMJHteoHpT
k/2BjRSHCoIPVmd6OGVu5fEcVw+U8/gUi8Rtwb/5kGrA42VQ1BoBeC+UFHVoRkyN
3Gq+8ZGXEX0ELWRTjmuTaPKkyUBKuFt7me22fwMz4BuZbHnr5Xh9azDcwn5WBRyH
LPAYgs22sZUMejIa2p3w2RNvpY4aguLzg152toUz/pSC0/V4NmuFn0IPaaLi1rzQ
nECVSQ2f2zA3oy57hQ8MkCSar77vhW1z54IjVBf4qVCjoH9GE1Y5W/qGKBTMdY+X
u8R8M2H3kZsd097eJKwnj2/RYDZpXVxgO55JWm03dgRviEQi5F6fFEKz0gEH1ZKq
ouG91DTxWaMxi4ZcbrfPPzF/QQqlSst9b1ej4iIPPxcxoGDtaE7fV4//1hAFQn76
dkMvBjcZlsmgyMbTAIW5Rdvh1F4Ehj1qrD39+PhJ04z8bQj6iYHmGQ5y7LR5ufVj
EGMsjICBqG4NUd9K/YSO9XYaR0Gs1zMVlMuDLgAnM79S9oAm3FYPoKqXuTbLBnj6
nkQ36OI42J/y9ujzyyXXgeuQ1lytWfgP2iXjnBHjLYrFv7YNdhNCatz1ZbgZ9V+L
sycQ/KqdVMTAvHLIgMRuwnFUPe9PajQD0qcQBPrj5esNcQKhzWhmqOYAW0U5qUOh
yh4nXq1CibErZ7QrOrgurxhyat1xCllnSE3gaoGDlkZnThuxTMIzBcm7nzMAUy0F
iDZqkemGsEjCf418vut1h2xxvhW9llTZdAAys6ti+2iv1TuaXl20p8YGUh8WYoFR
KIcSnrxPBs9Omo+10pxdtrWegS970c83t/83lRtX7N9xCCU/nuGMCMtwAm/XBB/0
v09HRametIf6LjQjhUQCYkY6n1u5lbhkOzD+WTtHVfJauf0f+s1qMlvqfvSIi2jy
bPFXEgl28Abj3RWduL9TQ3Vji5tRzPYsjif1QgS5y/heX3aygsNN6Gm82d59g0dA
UV+IMctYQ0VuQrEnbFmYsZRG0PkPw/M9wkkJGy1D8KEYjxUM0MmD/X0sLnduvaN+
t8DLgfPBBD9AMfGA+p1sbvBVVHz4HptKzBlkKMC3Q72yhUQzGgQ4GvvC4tQh2HXS
Z72TJKOnVzvw5PpraA/CieCGOrTdChXoD8sp8+rglJJPP83qgvW6L57Hq7nDzm94
mFkG81fItIAhhSKxaxMQP9Gv9u6dJSdS0eXf5HnMROAdT2q8PGyA50/uylynd4i8
SkLMB6Gz/nKv0qS9tseMQQ7qp9ctMcBNtEhsCpil/z+SOwgF2XEm65e+0wtdSWia
BmK1DMIgLWj1NsPZXWQIFny8xEJ7z1h8pO17AuMqzpexiIUqxuRlgeTxKkVbL5pp
/a4kccxk0Bzii/Rd03eezHhI1dKKolS+7r/Vn+47DG+xc+NmPl+qXfG4O4Y78l5r
ooeP1kIlaaxz9S+tHsi6PmKOK/qGYN4KRRn5FZiMM4HqzSO5oSMIPQ+YnBfmqKp5
lPR9wxUcDMKa/KfUdFKTH23GZjB6c9+xC8Jj2AhYdSX+L4UT1HwRQSsiyua78e53
X1BtlQ+/KZpGT2p75SV+wWMMyH5LSxN1aHSTpu/ENKbsYowrmvWItxJmFg/xQuW0
vrJziZ4cm02dlreOhUpvoiWagxufPw8tcJrgbLok0RkrI+Kr1LJWZWFq40yFg5tu
j1FRiGyZHGqu98Q29gtEl4X89QCGDSwQ+IqTLK882yXY4soHQSHCMvp1tPezT7fk
EE16/XYJ/42Blk/bItjyFRiZMygiDXs35pXI+u4RhKO+eXr9ruhCwFx1Utr8uAdE
r31iIjsRDHk5sXAWJp4oAnCt9Ab/635b+ocax+la3oS7FSwUnqDyqhkdk1XEMOna
6XO/zLOWv0w1ewC07L/IjzJa/ldkoNct17typfDMV9eh4xSDOz8STgdwrBWgu8Pw
BRDPatC51sEdxGOoEJWzkcfghFS9vMGNnWcCNKh8BFwitIktTpOkAG0q53rmHmr8
SLLVGplBl7COJKVmzGzxobJaVR7DfRKpvOQK1R6XJkXjry+l9+sTi17xMV5Utz3c
BKf2rn7huytXSRed8TvFIfyIuUi9ucLN9JErrD6OEyomHWhdSpBLCOU7KXBV0w+/
6+LG09JD11u1IXONrx9qG5Sk1RaBHdt4m9EFh1H9FwGDqjWB2yPgQQL2I4jhqK56
I5f7n0s4+X0Tj90ib1wDRWg7N3uUw1UUovJudOaY6fcQCFc2shmeC2kCdlAJjNFF
cKJLtAY1ZhJoQjDbBxln5Qg0UcH33gpRQYJjqqgQm1E6DP/8KwXPW/Ct6Ki9Mr5t
5dvVGIZE3dIw5bCPKHK7FdzcBsapOCESq6IT1ahwGCNUXDgjJF/O+0vUmwdK0IBM
08Tea9cYGDIJkXlvnjADWQQl2/L4d4c0LwFiSZCky3hjn1brKfY+QTzlyv1kuiXk
0dNqi4EFi4x1HJzxBYP1i/juRLSIpwknEiKg2A2JxnoP4wXk5kuqcrtaC6x/Bmr5
Al3HM0XI+nyQIurA3MtWaSdH2G6apWvboPo/O7gUkg2Yzqqc/ThrbGx21VZuzgnD
0kel4kskq5vZrboC0UZlrGAWDGw8fTH+qLY0Oy9ZLOHQm/mAtscyWFGBN2xnv0tH
MLndUSIK1bifl+EHnC8YddMJm5PRPJnYaCgZzPvQmXk6BWuWxAE2jDVx4nc1nU1t
/uVA6QbIJri22QkldwXv3B7sim/ENpbrgPTNrdZ+VKixm8jyhvHuEmPgDUjTwFGr
Kh3cjrjbUkThKqQpa1ue0YhtRCMSLXCU/bonj2PcEhZfh4mWkq3oxIYfOd43zuPE
vKSXNDH1Q2AXPcXvzUh/s0/vK2K896aH9soQRHkBucq7d/87e3WyiChN59V20xt/
l0tXZcq81aKK+NA5gTCRcp1ECmBADouJg5uYXJTRXZR0mT1ek1B2o1A3wTitaF0q
vLky7x0OOd0SXdgoWKws5e4x4DoH8o6rBeFjIAsAM3/93wqWJwjM3+THaJpR87H7
te8wFmIh/S54sZ7rHUa+i7Dnv8ZoemI08T7Fsdky22Iavxoevr31ZAQ8ky13FsyW
PTLgRXd+bwHKqRrhTfTtbgMks377bpFAzakFG68+U7mQ9XALHvbEPjtT/TzxAzpb
fsBQXKznnENZpIdTNQ7tqKUfuMsYj+CqHU9iFiI3VSY4l0NKhbBBjVgWTCF7EIG5
OlVnfBUNokizYTnuBRFUjagc7VKxMjFvL+o97n44mcFkpaKAD1ms24JlXK2VJsoq
sDw7zV1m7OG+9aLQHFw/dmRrcQD2rgwpPywUUS1ssSd/kD3F8i/DDy7C3JZ+6dXr
8UCcMtbkT+qSCScM6qgLekrf7KeAYIRzKaEpS0Z2BCxnmCTdlSSvtcoiDIK11LaC
ySkE3FYBHdVhzUN52Z0A2lyEd3iv3c+H1r8LDgP9WTRN/4djqYRMS1Ub9HNt/oo+
FC7UkLk61yPKMCQIbfnaRRCu/cfxVcfGe86ZfmbVkOwkyDmr4ck8KH8ggf5G8Tg+
oMCbJo165YDiUI5vVufqRM7R88a2i31dSId39bJi0M3E1Vz09HrwF5Rdcn02YgV3
LGF+8C6UmOdQvdAYyB7hEppOxaGtUTGJLNnxgb/SHndSeFJMguyinVp0+zrYZ8Mj
/AXaJpRjQ3pxOExuUhzOdGBgWDw3+4lDXQKJGf7kxK9vtRIItGXPPv2LmOwoD4+w
bdKNyLvM2vFdB3HNyfOTkq3gNNTTXDsmL+LINGyO6XQSA9cbw+s8RNzGT8p8R7TL
d+kM9AyXvmbfM62Iu/bVw50fyfAIxucuXK80+1rVCkQSWyc95UvAFfYtyEHfYsed
a26xIigV1/YqBC9OmlH6vqbFQPtFMWZDu+2C2Hts/RBNdGJ6BsN/4WTH1akLF+QM
3yoJmrWEQxllsc5hAZEyAIsdDcsJNsUGg2Cvk6OS60ZwLsacDRctdH0mhdvKHxhU
78o2jR7QMrJjD9oRssRGAtCS0UScn6Pwr2Av/PPrfa6+9IkN9ce908BHreSv2YcE
ETII5slJsYPZ/1/u/FGbqfQp1Hb7cSr5oarnR7HRJf+/GGF1VVB1oLIznFEa9xSr
/4lZL0MLh6BounjvdDEStf4aIsSbGVQavGxRLSN/MfY7YjQsULwvvJGq+Fpgz5PZ
l81iqfD55gh8/Lno933GyjIENtgX0i57IucXLLEBS41ZqardyyL0MT0ZaWENg5Zl
6uWrmdIwOuOzIl5UncP+5eHsd0994gqr20b1YhDhdKstQa7hr1ziiBGl0d8AIapL
iHplxGmZIBN2OGPd7OPf3oM1o00wJmal1AqtASlfLYypPSPGeQXOa0K9CpoJQEGW
lITRvklCwLnn6NXmP5QX87SyfBVpJDiIumTT8w2HRB2COAhCOHJpeXkIPa/jEFsc
wi0/p1MmfnXXcDrq69HesLAq8GS93cjffZbyRmlrkJtka8Ri5Wxd29agrA6s7IBo
hVDGMpRlChXIPWPmCTCMFlYqyh8YsaNuSvO32cnmkfQVtPYXKmRp2kmSRshiu3D4
yPe5F5PhxUH0kL9/otlUogRo1a7fgJ70AYGDxVyZci78MVEG5AvKO2d6urBeHxhP
a6bTQcsQabm0TT2WA/e0JPhQMleElczBP3ItEGNjgjsapG2gyLIQ+ExFgLIF+voq
v9724d9pFQotPl1jBtBVdAe9UkXJ55m0GAOUIF0fkzIw2FLDElMmKZrywIjhWXoD
BeD0hyJoiKwRmhMo6sY3Vc7eb7SpsH98LEHuiOsdzoV9AWs6o0t2NjfIYhKnQIvm
LopIrrCfECsPzer0cRcTLIejttu4ZklsfvUMS05tI2YeWJjbUHIIcKPuIn5J80iL
TFYJzO3czWb6T6dOxJ4Ywe87fnSOMXsf2XdDfI7qphWH1OFvEhhKABgY/RHApQS5
27PxTFlK6VneL5yQ3Xfhc3yrnmc85ZO81QtLDTcyVwT9DqWL9p2PQD61si1Nf+3u
i1iV3e4nWvFRZAAAvHhqqxy66qGa06O90Oa4ZsadbagQWiFZLRWQY7vuv/5GHKZa
xhhGv/w8qSt06SjSYuadRfyoeDka9KL453y5814tZYWSjFAPPol6W3WnJTSO10r3
pspQc7eCXiU/3NYHywva1FQCCNv4tMIQuFfyGQiCgB4X/+VB4QxsVUar7LwwxlgT
wEqkgFUuF7V4oZXjvSxQnelkVsPozmr8NXBB7id41zktBvkUggY+IogMHOPTz7tA
8pxzDQibjIM4WZW7TMTAj0SR54obTx+H839cGBSoJ3s1whfJ3k+836lfCjVzSscE
a/FmDgcRpL67D2++nrE34/dydQtaAdBfLWKKppUrJDaveo/7mXnwCTwSwNiSQh/Z
kkhCD4Fh4MfY40DnI0eNmuD2F11EKnPh6rJwS/a2YvCjV8b9i7KWiPp2SnP0cp5I
RKQjcjBUluozu2dAKaYVhLuAImEZX6fd1cJEApFo73lCk0zF4F5vgwOqjvXba7G9
XiMpfYX+J51i+f6MUVWIoH9zdMpUTTwyt5Ept8qhLZsdzJwLJRMThtJKYJKlmqug
8waXkaZl+zlh8+7dIXp30KFnmGrwtlvNWWNumeA9qSO0+PuSyz23Kt1ozCfZztcP
GzMe/N7Z0+mfTWlhZUrKQU8CymBiEgeTJNvZ7Osku4Zp0fGKHY09I8RhTKmRQe5k
hKmflC48txJsp8ObpTmjNWgGXngsU9+yHpg263z2WKAX4dJ9jWPHnCbkIW1xbNFY
PYqEokM985DKbVexMMQZ2qYsd0mPlQ/k+0c+mAsVXD4BWeXHmbqnFfrkNHWiJ1ZM
bsW7XROcwV/EmeEpP4DUPPT3vKUczM/tmRwzdgYQsQF2ViNX1zghmucNmhvVtOlP
lrmHufq1Mn07OA68YRgs3j3xkTzpYwq5DjsGVaWsEu3hq5/QzJFFhhPW4YYwRIKy
kaxNnZNvGsZl1SS5Bnl7Js4E5AUntH9IJtggk9iTs1QTCC6mCzcGh8t4scZtT9iN
OkKTtFwhud4Ky7sKG7e3U1cwFar1YAH9ee0xw8Plx/NJPplOPTGTCoKITqhvpSlH
bPsmR499/8XWScSwaWpbcVb53AmT7uL98Nl5U6tPDk5TJ6B9Vi1ek1s3dUAI+pJA
OFa41ywfIuAzOnsLRsAvmASt3ByLkiCnYU6ErWHX5yNz+IuOIulC1vBR7N3Ir/7B
ytOQ9pdPO+Ho9Boy29Mv+KKHbVQGrpPs1ERTzqwIuylt0QWhq+2jBiTrNLti8tsl
PfM5Zex+m1JPk9D2DKw76UxrG01AFmYx8s2tE3yBsDttCw3OI5tw7ZFm0ZhWRFsx
8TJuAgKDHP0iffHuOJYjuN1BZroRbWi+qJxBxk/KiHf15sooK8CM8oUciXlnCANd
C2e8puOtYAZV7Gw7XO8cFSGP4xaVnBLSTjKIi19six6busHtqzZDpcDILxU4KKzd
9f8e2BvtwoYX2+0Alld38Yw+sjWgUYZNOXimXZGLdVvdmMLSm+fz1Q10m2H/gPRJ
he8CnW5fGaA2GO6uChd3/iGcUzO48y5EfCIiKNLGxoPupdCzppB8vi620TZ4N+sa
VGPvo/6fLC6lY0fP+Y9vy7upKT6gvRQQW8X6CzCb9BJjrOG05vuMUGPf94yJuG1x
MFxaaZvFSPGe/7KKToO6YMK977evKEbGrMzJ7zDjE96Yl2nr+V/OYj76mCl74e0I
BxaGMhCRXYjmK5sBqJfUK3+IgBvN9tLSRDw+0bse7EyjlXqYI/0yQ8SlNWPRSQ2z
YoXjuK38M4WVqq2UjfRb5ptPvSXy53AaRngt3QkaqtJJSPcuJb+X/h8yqjHrxUz9
JcsA7x9Rnmh60hsaYGZdRyljbuESKvtgObT4iT0TqGqefa1jIuWUVuPAfgc+DDB9
EZbHpTrMRRFtZLVCkBRNjy5EZfAwj/jfNEeapYULdFlY97TlqwkbCn5nFtqEPko+
0gIn9dtvs80Ucqd8t4LW246NgKSLRgLabLo4AefKzlnVp6VG1iJq8Q+f3vW0FIzj
Hdrf7iqwWZ9wvLf2kFOyQ+VomSyGDidytWiWzAprEu3hAHaREJOy8OUJ1dkwQ1ET
QLnfbzPJXxIjjWQEf5dt6Dthhp7FUr+9kaPoMGbZHKuJN0tBPxooBhkI2hgLXYkp
aC0NE9wl0rbEQg3y1t5/eObugoHi+t0oY8aqojs5gtXvW7Hn7kLJdiLtp9f8uaDZ
LNjHln9cGamLVNm2ODccUCDU+PQTymZShvUVI8Op6LbAHSpA4hDYaHO3M6w7Hs6q
AUo1AbmIz1quU8nKAddnyGNjlojPjpI0y3d9BlSyUH02VKHgxo0HXKXl9qZS2Rw8
nmYCB3mgywc28RX9Kyot9XHJ+RjdRPBpFra2bta+DFvuL2/a1aY/1soS1ZoKGdsl
8n2XjYzs/863og36Yag0hNZoYmnqscFepNR7BaX2jMWZ0Bga0JhE+avgC/VrV4wv
F+kkzo/2PjEQpSxT9JIFoYs/+FRzhNv/VvSNZ6Cja0Mm/xikarHe/B324MHBNluF
yBzxjNEb39uST1Hx0FcOckUaFrGuTZgp6zfiXtSOAzFB3c0MHVPOzPJTh+/chJ4b
vABeaoM3zs6fUJEJbzFpcvA84g80supTSXH4hSWgXX+8/N/gKR+wXdBCVq2pIlMM
bHb9FEZ47FmZKHSh5fN9vx/iih6OFy+GneqsaaB3nLY3ycT8SsKRDQaG5gQQXOTI
Fgubj4PNdNPlTF3IzoJPGiH4GJ+Xl+CNh0yELIWglG/ArRvp+hzdhF0keiXUiTeV
iujJfgN6yeIdwlzFudjC304IZHTjK76YI/CyRL+m9F+wy11PjD3ejSB/aSL/6nIV
Fl/sEOFOggzqJBK82TCuJDyn4aQZP9b71SlSkFJfTzbngMibziHCg0bJFWnwY07/
vv0xGak/a4i8CoQbrd8tOQlVhaToKVFXCm1mx0FgnkLvWBEDFQsuzikQ8gDa7/aQ
w73jAT02kx/1ALyo0ckgS/yA2ZAfzTPAFztWZS8exfHaJez0yM0PEo/PLTdkasw5
ChxCynfwqkpYxaFO2QpvmA0ZhVa6PIrC0/WFXms6PML1xsu8Yq8GnQGLYxZxurqP
TaITlGfb1dLT6z6YcnqMjN+04O8l96fn7S8YejQXvk3b7vTGqik3tOEPAiPRIEv8
arZxEFeJwAoXHwRlbbbPaD3vauHxnlHZQBykqdiFwAgU19iR24jQWR9yhdbts89B
m8kr6+Tz0zRVOFitlKWldVgcYu8EcBWD3VezJhPI1WkXG9AEARRLHhVFxMUXJUIP
CIesjiWXmOHvPPwVejFJavF5vyn2unZOa986GkFEz7dCCSgFhdrdcWdmSv6k5WHJ
mwa3UUOecVZC7PSGgzSw24Lvp9cuDLDOgR4B3smr8+H9BHoyPv6ayz/LPs5eITni
u365b4bPhlKt+guwlVFefIQy8SxeA1c+e4szkuBoVjV/szi2I6YitZwrihDfIG3E
XfOEvfQk43auoECqvtq2OqyJ1abBg3Laj2tWYbarK80fO/eVe56C4jKodtdGS5mg
PJU9KrXDrIG1jZ8kOGJGrNeqTKX+3jimIIU0e1xnLdmUGHvJioNstUZhoy/v96K6
Eilil6U4T0Mwi8jQLoqlcLQ4ryEGDBXhuF4OM093MFVvVfrZEF+A4FDIy+qbS5sr
7RJ/uFp+W9MTJ/W/QXoY+sbTcs2Riu3xLFduJId1TwHep1WRzEHyTqnyd4MmgwZ/
qYkErntq8q2QM8a7//4SghJm1pE0u+K6KzyzHhRlrreakS1vrLP/Ln6Mx+84GXHx
OTCgZpn6Ll7hKgZ5QqnXBaMhA1LBnpzixZwau49AwOtswDdIHo20nifm+gyFUvgU
EmimkYzie3MnDqumHtEDpfoFPIPM+db0VhvKXcEvJeclkHNz93bOtPGDeFMqsbuG
HFUQr9joOmSIFNZKVI3ces/x5wCpxX7qzr9CROPk3AWfWptUnQWC/Ob3Sr2ClyCO
XD02sga3pdpPSo0DeFu7K1PqoXE8YQu3oD7PSTmjCoTHPwu8b4v+aujH/ZO5EViQ
bzTK1RRzxGpYFVHFrJUs8Ibvf5nCOHmnVd8vWnHNlI5DL6/WrQVnuDHCiHoPbmxs
vHpMd5f/AgrKd8lcrSQFueEfl7VbUEr0sMqylHABbrS0BjlhXtyHvWuoYC5v4KaM
6ES+EEORlUOj2hViBJDffJfHzril5R2OgpkhiM+Xi9jiIgTkUTuE46+dYzJDbKXN
z1Ju5KlgX0v/NBQFpzr1xaQ9oBxa3N8Xph54H3MJCNrPo7ypyJEGrMLV2qsXG18G
frZ1/mUrySJ4k/Ig09sH8VieorFSkbCE8FytX3RD/SRs7WPtlLYhXob5jw9LUY7j
22vrPSsAMGTBKhZ0eLXYKIC+2idyGo5vKZBTOCSJfLoN51TQQzSI2YTXeVuStJwA
qKTIzQ4bOr6KAA4uju5gD6KxNr67LpAacaNgmB8IhIqG6lIBShiacLf2jZufx3TX
SFbwms06XUpN1QCv5xXkokrDG1P147H43V9EifZjq+Jrv2Yh4PBSMoRkAzE9EUNI
47nFPgFz23+qII5/MCtx6U+Ry2bDT9MjP3h6a/lFjh1PSeBjxuLMlqPOcQT/PVfy
c227dH5qkpzDBwE1RSE4EP6DMcvj6fyVjSByEBwdbcz/liL5xhFxNlw2+z6Zaiup
t6Aw+U0Z/8BVblwYSr9ku6MZIsKmVQvKvrSpSbb23CQgDpzwRGXwoJa7ThZSsfea
GuwtkSdF6PpEFVUv6Ag26dVFbc3eIEvKopa2mQGAiYfweWaoHgJMPXS4Gb0xDcQF
Ye7v3Z7FTCFVNTH1+nz2SEWG1o3mrS0pbe+Ao22K8YyCvmr/TOdQSLPn1Tx1W1E7
qCB5Zv9R++niUWWcYsqgTkkJ+63tjnzK54iAkUCx1lP09GuUsl5qiXlYC8+tiNMG
S975h9JiZUaXA/QRzo3tpSA28L8sa0t5W1C1mHniU5VPLrk3UGmvQbBSzpueVtAy
DjmpxTSHsMJ4PKHQ3nOgYjUnE0A7PxNZmUnffkOmeFdxOcR7AMrKZZq98JUfYt+f
b9xLdijrphnT4gone/WUMW8yDZT4I/NjbeIrkCiSj0+DUxxFQ9cF7EF/SvhBPvYq
w1EJMzqsNMoyL26K8b9a+kOdDeGu1TKo1sWu3FNS+eiRjSvg9crzsqPEhzYeTfqV
2meJC++GKQm7n9WzcSiXXoQ1NLLNV/dqCP0CTazpapVFOYm092eJmpJojIY0klpj
2dyvcZYIaeAvBc5PFf8ElNkPh6Er99FJL3ysyyNUrEhYxrI3R+KWHSGNYXCBO+Jg
OqEvcrvZl594SpKZkdfuwys/rmVjJSBsCFqBMtsTMDHhbrHUFuWLMFn00JCXoraQ
MdMdlUILhliI0eULHZXLl8btmaHlhgvKQMK1NV4dqksFtQqh+PNwqrTUMMQ3vzJf
aFVbIxq4Yp6WL2KeW9spZuUKCnSHg4yu80gXBXmN1AGIAEMpWf12BffBgMXyNeHi
FqH5961QpPaotF/blQZ53+SHU1/1pVCA0N1ytw9aRHLLW3BuhBWZHzCnMM2FTSz+
Y+BAII+hngVJsM0ivI4BXlvb45Stte+U7Bgndkg9oYp3Y2gO9ID3PRNze6PlC0pp
Rqgq1C0aIalbBq5Ely5LX1xBl8dcq6QIHqM05z2hfbhSI7SNvvM5wAiLK0Eg3Grl
06Z6iEsGacGq2lHtw22vL5fYFeC6n8z0hYDawh2IBa1GbPz8NQzc+96u9WSc5aqy
eLvIjtfPten7CNEZntgv60dex5Gw9qzmGddL7dbtNzdfE53Nd5PRbHxwL1ibfFs9
9f6mJ9lvqJx9Fq4su4kluii8ucQrBUhxP3e3koGFAAg8be4xaAVUVxgLnXKkxGTI
VPX1WKwNcN/qEsDDqdMTyX3UGfplNagVN7H3wUtrxBFbBX2AV2szz3iWvfXPJyzh
z7p0VAz9OaAJUBIgpVXVzZO59fQhi52tu8YxvPZInjGYg/FIYMtP9EMVtO8Q5LHT
4xd4yldeF22Xw5XjzAAX8q/tOC/WAxacSnY6E3lmff89IXlpMKCUU+fHFzntkyTf
+NkdsNN3Q9i3G9v6cKcMIkYyoR3Pwef4u3itqO3sbFWuCtRHprvGz8+/Ieo54hI7
8NfhhmWoQXElOA7Sccf8BDZ3YA6bJnE5+uyiVNK/f50mMDZ5CbGIhIIHqy/cnAQG
iX+15KZy5D9NMFK5dynz0AidEyHJqmq4QgK4naxB1pMYnGHDYoPJ8G0jdUscxzu9
H6FWI85t+v4zkGYaxVu+zau+DG+GU0k7wX1LF4nTsjgw0pVd4Oh0Mvd7vFmOWp1N
c3LmiiYf6yVSjhH3RnwlSnVsEuPnG6eyXTLitwjXQw70lUAEeWgPCqGG9O+LDmj+
b6XZ0ntZ32YJhLsZnhO7YWD/294edsAeDmgmgskJ8zpp8L4TKnVwh6bLThU2qVZ3
iSe0V8QljczNRWkLlC5KOA5x1/RDfvHUqNKiTm2yBaf3CC4ns4FL/+WBh+JOxi7z
WX5YglwF6Wzq/wVlSBkTdgAZAuthud2w3lWghSbfoatJJPWUHX6y2BJ2d7DXVn95
WtMmzsdKxnO7ZD5mBxqCoWso5dGEBt6SEgeCGM4a5VVODmqa7Bnu4M+nUkSQ/7ze
R5STnPVyLREV/JFmdqoZxdZ0TKAKFVcFDf8TBaQXuc+DsfnRvwqe3JyzPpVhDoGI
ckjPOIgJZj42vYnGAlCUp49My5yeLW4E7Uuu+ivFM5B7bmqO1telbHyiVxCIhgVT
Y0CJu9hl4b6idp3ELgT8zEi6ybw/u2VTYFvCCv6Lz14tN+prbYUuslWMyVhbLQBu
bwA5RJpz2TZ1tOeu56/BtjktqrnFXZttY52OcxB8oMVr2Id73+Vrw+Rjv26echiH
akU8y/n6++97n2LAx+9L6TFpHXgn8+26k+q1kdyCgpp7ETRh0eqWLtMrFambjcSI
rdbtEee+Iy5gkq4q6Ae1ALCrknsOmtL1WUaLkLx2xaTTo0ScD6hyzn/LGTcjQvUv
JOVCoHI0+xOt4kAZdu7hDDHkfuorT5Nbr/UzBsyItMjWKDagIqMZvpBGqC2/cYNZ
spe4yfXZV3ZZ1Oi7IugIBA7+b8KyQV3gRqKi6dkDMasgjsldUUO07vrvG8AnotvH
2AkPJ52gA5uGUsQ1s07R6Vh9AbYn31D4irU4E9DjbKWvaZ/UXd+bZ/7Zp2TDKWrP
2ASOY87NCLPYA06KEs3qrlU9F0nt7nIUfbSuRfKkqvyNe/E/6pIf/F/oxxCUtkXJ
vWVPL/YzyK5MGIs3gssO0dav7QZHJnF0vji5yCihX3nZlBbhD0npt1J6ee5df+WT
kOtbhJ0A9SdD4pNteQagiBR/SBaxCtQ4EmFrGh2Y/CjeemWIqFC1cC77umpzppU4
yVkOCgYz4hM3JIzHKvY6xOUD8aojm/EXXFOs4KLagCXZdN3amyQBiIsw5Pxb1mZI
Ljd0jrWzQJg/e9NrQwbz2wrFEG55F22zn2u9EPLMLb1il+k4Fv5MIa2/+rpmLOCx
DOqRewhdN93WTGdH2zSz0WETkRx3k8SWglpIy4avk6Aq1aCM4iOzZ98YBQn5Hw2u
Xl4TJ279H3+2aE2PXfq2xZhWvsmDDVx1hCaP7FVgKXGnLDHFuqy5MMPjTOcjLuOm
Wczt8v2CSq8yhQRCM0/iL1KnJMAXfijs0jgTsi2vbAYiFdzrf38ji3EeK25b1dL3
xiu8X+fwHENdDi3+jrGrOMyI4uM9eujQL8821gaewvSg28yCsCzTT1lEUywTxK8H
Xk5W0ivpfuCkrUTmotMCSbf6MX0NF+RVTqXFxb1ItXAqd+h4ou48+BrA01S9CIjj
aZj/IDTaAEt0lK7wR1VEdF00Y9Geluv4fUY38UB/vxY8vA+JUSrpt+lALGv3lGPz
OUu7kTJ7ySokMQmYsojmqDoS8X0hHpWDQUJPGwqGf6KdVGWqiP13XUYooruwfzwG
OMpmNHun0LiuB332LAE0LNbDK1VJ9T6mLrcD+Jt6ww23ljMiUydo5G9cpVg1Lj9m
7y1gcqGT5M0lNR2PzYiuiyJkvIkxUmmy/g5dRQD1SrZcXIt8yvHd4LcIj/LNPtXM
VR3ASEBPTexAjXmcfyjV1Adz2KWU38rwVWERbkpJiwXbgfu9USVTPl6C9pRRfAaZ
EaQLdqz/6bRw4HAIzgmi6Qlj6ukiCzrCSSdsBO+aXvpGUQ/wKMu8uxFTigYBt7Jo
yNsW2Gvj6r/CyCB047FkS36cR1DE/lMKsoWG0GCtknueQMItQdZrlg027sTX4sIi
0RiuKXvTB9+q1PMDiAI0pW6oLsYyTZr2fjlWIbrJZAhuP/+gHbivO5+blUQU4D9F
xFwBy9ucaZH6hqSnG7r7EvtEjTbWG6QQAyp7pqKjIAWnqBpVbhyAcnzlk+fSzOH6
3TSIxBN4sob5b6guDK8GQesn8Odsjtds2hP7OfP18BSrOc1As/SCSYLG1J30yg1n
cjcP3JBGKcKG2NLgaDoFMisEtI6KrBGzDYaaZCEgi8VFKj7bWiEBRxrwkbVcYaDa
fJAvK8a3biGMLOsBl5LAMhgX5GvG2hAEZiXG2c73u21EuQW4XLCe+TsH8bvdfR4M
6tFc+Xc4/XQ3fF78bl72AA6oviiMcJDrxDAt0uX8Z8mzjk6M/eiT8Hb0byRPbto6
1gJMUGk1xn831U0b5adtV9IMjQ8d4vh1fm+gtw6Y3+zY8qFX6/u6dAkHIxFgaw29
Ji3HQJyZamNzq0Of5fs6cSA5X0r9KdqFLhEYqqsNc10ETSgERdYGaJluVsVaLAJU
iT6don2uPVgE5BpKs5CKhbBZHTgjZcfExEpVbaVwnw4/vI6IpFe+1PaoQT3YfbNS
Z27bWD0+lYOsn6c3CQ42/1I6tJ3KG1U5vQ75nYBgR5b81L1BIvXjKv34cw0rxZdb
5feCobDdgzvPsqKivH12didJmctEcAlihQ9owtAfd61d28ZAyTK2oef4Mc65dUDu
S/zpcRY8yk92kbdG7qcAOMym3PJY6R8LQkkNeR4o1WdFsFipppYoh8FwdWqXQQkb
dZVlWTVL00JMWbO1nBzUhe8cdl3tp4hj3HNaq5XkEpMOwBO3fJuXIm745zD7/5ro
ecTP+wHV2OXS+DtW1ZVRzbbOlFqeQUTFT5eRDbUdNrmo/gkl4pLU3sF1qhUkCr0+
+MF1zvLav/H970clZSoWBGJFF47J61NjP6UrR17LBSlOrfqFq9HdZSwSZO5+PVcd
UqmqMTdHMGuhCHuJLojTJ64dOVy/7aI1TQliTeIOjLEAmX/YvXTpJIoRXmPEz9Ed
yydGD/anwweWJMkWkBjBvzMBblbLvGNO6ADchcWCiynNs6HJ7F0QZNELSgqd0BWq
GFCEzqXA0v3q2gwHMKrXpAhu20U028zPJ3sShlkWM0A13yqAE1AO5A9dinWs1rSa
coadGInYrWv3lyPY8Uiu1gCFAXSiRnlPYHkz521RFbVMkIaM8NtTT/9y36Dh4xVs
FeJ8rvDxtPBd0I+FjyaWy5UzkM+X8a+GsHfcqCUQkEPWtU2RAqgvWhBzdLImxCZG
4OL+LBCPUp7BmAdezz9/Y4gZJLr/uinndqdlr7IOV8AwjppUaJ0Uj1tx8Rs8kVKl
wD8cW2ZPbeeWW4ubl1vqkXQeybkoeuqSIUJ5TNCKspIsCILFD0vXhJmVKQT7UX9B
yRvLFJqfPiNpBhGGpNylgq35BjopdQ+E22KOOLeTZum7smAMY40qd7yEMPHTdxXq
0TPY7ItEuT8fOFbdvpwxpBxpHgGACseATOnM4ozdiYOTZ3bHderpg/9jXHeAfv4a
5hEkplBzO3lxpUo3jOJgOZCF5Do2NEH3S1C83v3xHAl9RWUkwX8mFfESVo2ZOgfr
QNBbU4rCwv/AC6pz+G1QKuM17iMqWGMygsLyPLrb0sSuD4zaXRoSzA9/Wx1ZXyzt
MQyNYBXxyPIYKfea6y6wlFyXy0o2MHSfmmf2fmNNoVTrE65lcgsMB7wt+Vp0Ovon
m7f8KqvGTJ56l6yW4D4mvgLT+P6gjcLh/02UIOT5xL2lVgCdB1ruFdUstQP/WZhH
CcWkByXElrcFcYi/nvpMsGMuodhD7vbndcNGazvyGEaoCsgQRntGLl+8NJrDeFEl
kagomXanIEoDspu5AXmFAUfj68WNFdlLepq5wcGUJiMr1X51jFU3vyIpscNDCLgj
h8ScTH9ybiUnAJAr9UURqX/H+yHzbjM/RqMdvGnbcxj27eal9k63gRpukF5W85Bi
pltV3cmotFaJ23j1Q9gF6UrwCyPdRExQs7NecjsetUWV39xQekBgzXR2zSIZDcNw
b7K9jUr1Tq73/Ncd+oYHM3r3OgFHLzB9BtCAsdOHtRooUwvI4LN6U6VLdPBS0FqX
ue3CI1Y6HLFSSK61cCfOHFyGS+FpPxqA1AvBPoZVp8rbvGbnWIKCyxGO4vg1f+/V
QpOYV3+zvr67qgJ2gUQxaGdXnB0ImD8wORUIZEc18bM/H/Z8KCb5cT9g8mVEet+7
mxgNhxe1SD+cI9fFjKSIqK62CK4NdJxAsRhipTvUoQW9qCg9qjTdfVVNUs1rdanQ
mUW7EtHiLhX4rYpLCA8elqD2sFuKKbZP9qdNLANl3cm1N5f+swd9kdsPLR8LjpQh
v//sn7E+vfTXpn7VSn2Fh34GbBxsVlJ29CvRioHu7OTx6nd65/qXWYBMDclbjzBJ
ifOmtKPFy6s44s+L1qQAu/pJ7ZEijf9NCkSRdeY5Rl+7wNltGsm3gNYKTgfstKxK
477wlfrStMniq92xRSxLHaehWhAjOqaKoTbHHOQxvitzwJ35KvZ4LuPsUS5Y1Pps
024U+O++m6/yZbjougGR+XMKp8xcC5WsvP0zhCCNoK+959RUBOL9bNIGspD+mUW8
wptWoP8mAd1S072xzDp3/FS1xWIi0rxB+fL+3DYAm4Rsurb1419xoecLUjDUnhw1
KOGzMLBzELs74DtG3uKPOu+dxWPqT90yqFFGlIi1o3o3jfdfqB8L1YO2renWlMRE
45oi2PAMLJ+vBdzMAryzG8wRO/ql8MJYAbjoRYBRbqlyOelifXVpypky/wGex4FX
+2rUJ9ggqBcLy09+WQgMQGmj5XAhlYrW0q9b9Nxh3Bin7bxEaM1PhshiF5hfmhGd
LgHOET9bcRNcfIcM07SRIckHM/HeZlzLrITbhKLJ41megRkuurMAKw4cn8VuL0j0
X2ZxAVbTrIuLwtqNITPqhC9dfFQ22ld4a6BA1FRtXPRL3lAWJLD1S6adnqxJfGYF
FKT+0cwjsOOHfFtyDk6a4WyBe4vOTYJIu4d9ZaRwRiFFoE3dfMfhF4TP/dMwXHPU
J8YVpE/LuegcC4BNovoIhHeRFGPE6MV3OnrYV6YERPX4U6o9ndMPjxr+pT7PFDJY
24ogKc3wtwi3dQF72kVe58bix3XxAh7H+RtNruTiHeUB5c1oLVlcjqhN4E5hSERB
xYMxmCITlKyqzlEmZ/2c+66+RbOaIPNVO9ravnjqr86VU9AW/oHAn2TEPilXtg2i
VO9VIIkIe2MEIALvvaBvhxodswpg1fFYQYsEchgA/V+f/wsblYB18Eh3EL1uRBPH
q/9ubGoJFrxgHIEeBeWaq/Lyn0zCWkkzVhJKNScDyGYQGPmvHJfR36SWa4QCHDgl
J47a2L+N6VdqFfaBSTeM6nJeW4E74wz3w25y5bmMActehUvWfvpUUve737AP+l7J
gNZuIDXsNTeYBuUWGKEhn59/XxMy8tuM/Z9c8TVe41v9DS3vA2/OPsxvtVgaqtoX
deVCzog1taxGXF5Kx0n7BPNMpKUvIwKmMosXoRuXZzCx+capXogNpCgNX0VGfYVw
qVPTBSsZmNcFPt6392/UTHZRslJFLJo5A0BXkiWizOagAMXaTWdqBcDDi0ywM6/i
F0x4iWtOHV06GCN8YJvyG6vCB5RyF9jGSoxjI1r4xnw514VsIfPwUfeVh5WYtOpN
O2OtfHDdPsW3sWyYDB14AC9toyxl61i7s9wb5emBrYqFkczX6ayV2NO6DjvzjdzS
yQXTXn5oXWS1K/gHwvoUGGohBO2ZWc7/NbBHWnCKYjLALzlxocLbqd5+PyMrkfo2
oFRAPJd3aRGrfh9IgVlpM6tuTOliuSru5+1QPEshKrinWAoNc+lhWCL8LDvEyiwG
yB+arJJ9MGKWVjQYaRo7Mh4d/ZfSxIO4UGOZmZn+MYUMGQOKt9lRWIQ9Oxc6ssql
4ZeBaTA+8T8RE+hWa78c8T9iUWECYjwAtfYN8K57hJ7DKDX5StdRMmdC4k39Zvdy
jerzO/nuuMahb2y0AsZxe3ySAIKFp5PDxr+meSjMJ8i5qwpAqyZErpp5QiX4aeqc
4niCDG93+wViaMbsTNMqsb15lhJ9K5ugd7Kg78Zt9pkVVUOWBThbXBicXDiyY4ju
pMi+KLV6y/00TibkhUCFtTyXE37Xuth1QpTnhznOfihD/acUthOaNmg3kpP7PoTF
Dm2R6oV0/zZGcUAFxS6JE4HxX30+CcHsdinK+QTZRE9Y6IfBZwFIVOZY+u1MUWnu
vn9MLpZ7FboXdfj0DmsJ7kQ4ZlkG2n16c8KguIw/288gw11dTBxCo6493winMRTB
XeBCBMrIEQh2OdPeJz6vFMsSqCVtwBAflnKFzeIT8LqPphFpvr0WImXTz4iCe1vp
9rsfBUlss/tQf9AFMYpzoqwWOPc/mrRbhsPbhTD1Ftd0XUplN2IhMhPCV2OR/IML
FKx0LklbvdPZ1G0VEFmWHoSv5PVkBt2rLBewfRnkTLHHKQfrkZbCKd0TshC12T77
+2kafqJeLrCX51NGwrV1/mCgI/kEJ/n0iEcd7jroou2ORBDSxs11ObCzVcvf46/J
qAEdR0Fr5EVSERH99QQUO2i/aM5ZZLfQHy8Hbghg0LIH20Q0X8VTmGzRiC9x8UZn
a8aqFBEv9ZrcowqwQJ5zMJF463TRw9lyBezP0ZncGsa594R9KRawWvcUsb/GUrtF
MshX3R8uhlkwNh7+nvaEVXlbNlqhyL1O4zpte/Cs0FITUJotVFe+EesGSuT/RpSx
2iLQRdBCezrEwkT50NNgXrJSLUP5uN1KWChKSZ/WZGcgJrDZJkbEZx2wTKcexfUe
lJb7WRNUkO5XuTS2S/FmumYlsZn84t567pVH9PwZfU8xjM/pxHd4980/LeCCdm4c
aYj4lfYmxoy0cTjuoIXHwpLGL2UJX+xy6ZMjQwwkS1YDQbwPXuu0Tc4+davjNUI7
2bZC1itHJdXiZNjDRasI5qXiSYapL+NvxXnVznnqdXt+5GAgu5vmPKUbHOCtwwsC
jv/99RkPNUgo4sm5Nw5DkEvHGRTQf2APkamrQblYX+G+rMaFKvhSuVFUXIYEM1cj
XpvroYQOKyM2v1Eib7r/7CwbASdJhijVPS+P5eTBfIH/vFggMRiENDnuegNNJASk
uyXgDfaJBF/mqsNkBk7xqR4h/ITMfCuaf0jjsNVPGZj89+gfHavcLhdizpPQuHzR
nl6Vws/NEHOLz0euBPzvhI0lI/v+wBG9UUWIp33XOtjpJ7qFIbqmroouRTxt4z8+
0zok7mTeZLIdykRjzI/652GBXcixOewVEcHQHPN+fQ0BZTnPdmPWktYugus8oTtf
3peSh9nAP+h+Jow6HFlb8XD/2ww74EwsZsc3lp71VW4BGjtex2Zt7fxcw/l2Xqgt
P+x28oJALae/ReAQkLAOfVbm928AN5jaB80cc4wXP86DMP8fbyMEct4GT4ZaUHXG
E99saMX+zQ233aKFLL+FiM+UYxwbL9GQ7IvtrNiWh51kDEF3MLpMNBlCyLSL/wYX
rC3rWQ37kZZX75EAXPTmQ1ZT2WkXXgveyFhpFWiH6x5qBTvGgo599fhzyGLsaRmK
zj26eFCQN9aJGXUC3HBpcWHSb8tzQbmG/8MTcmhyKp45rYMO3BN5SGSzYQn8ubpV
5DqZweDE5rxE7WPKAMlP8M4UEq2B+dBmt3ckIowaotEavwkRbSh+iwEBpAI0SpbE
boWJtJ4wrtV/TY/gfkCSyTX6/PHiR/xVwyKq/yVtUQbprsPqBm+A43+TMrO7dhn2
PWKF698rEW575BJeMBy5ZeIGcIdPdN7sBjETLmaT/BPxtSETvEQjUVb03IOIthlb
Ig3q5mB3+RlCWmegtvHbG1ZH2A2NdoEmJQmJbfpPa78UgznrgjXODH1PpjxTQ9ud
0zqgOEBAXipx9VBeM62W7kWxtpTMbsyfWZr16oUxnyfOdn4P9IR0suBE2S9WZQIC
O9La72wUJOMKSxflkeyQ34huc1zzBckTPMhjAQaM5QIBvE+ztHBZm78Vql/66qi/
b2RBjSsvn4sn+ZQBZ9iaVhkca99qweeTjkRZj0k4cRK9i6Rlb+9o3G80f98DXh8c
zFQIIkkmgT3i6PvWUk6cxuLayD5L1YC6/kbnGmmqBpKbJeu9mRlXXzkfnv6P6fBb
saOaQheMvRM436qqKUOwmyAe4zMjIjYYYgrcdc40aj0viytrpbX0yEZOSBULHhHl
Ge+NXPKgFosOjh1Fzww3EeUCN8eS11N0scoKf5Eu7O8d/UGNe7ft52IqW9g42vak
upaIMXk3CTEu8Xb1kc3e50ffOinm8RxJx3rMwaItr0cav8o1Jigde7H8kZcYeGhy
x06dUTDQwmkwB04e6pOREsdd0ZogGHe2WCrYFAfUEv3kSHk1mPNF+JHYT98GRg3O
TSuCF8+im0UfGxNktYMgkQuMdov6a3gG0o6jp3BP1J21G2b9WBzai2AuCXxsCfgM
1Vsgagj4EKcP2f76fsowSr6wU2NYyN/5Fp+3/XLmYIdFOyGUjVuGHW/qMlZONI2B
cG9xf9vjlvCTOlWWJZSdBaHi1CcTdapJzw/fogLBq2aSRbtihRr9sdUQ408mjerM
ueKDWg+piFm7t3+LpWoiCgbf9+wgianKFl0OwQq+pnZM03CIJ4pzB3Xmz3p8wQnH
ughsSdhqDQ8TF44ZFXoXiQi1Xv23WdIR+eWB4rK/P99O7Rd5r4UZH2PHHBrqireB
EigZUhPddklkG39mPRwxfoNMsR4XlIq15MdXM6IR5E8bsRvA6zZLrxM1UnThNhQW
Luk57QPgMybwJIbyd9gC3hieQSWEloVskOrerSJUwpU8Bj8+A0hQef1lKLzM4Osd
/LaERGd6mf8OVDs3/8/BcmVBSU9JU32b+qSQCSr9O52jVVNmqx7pEDE7r2HF/iKD
Id/vNi922Lgx7Gms4B0yk5Py2b/d4MsmmKq5RnV949CCHvmS9Cffnbc+hPpbNKbl
GxfT/2h+U9xDhBIQzqQkHPLt0oQZ/JFIntteQ6EnCwQhkXfVEM/wqF3l3IrtZcWK
IJQxrIMZlflX33oxW9lU7jM6F9BZC+ZsFVTVbxdzo8/uuWW3We3GNRdl4ScJwHeG
AiCIUXrXxwhuaL8uA7fzoNTStnd4VBxxnW0XCeVky52FqtGbRFLKLPUA/XhJtHYz
jHhnJ1KYKxVq2/CMiOOAk/TL50Ol7hWS0HunGMUPxF3jdFeJ4lAZYH/YVsHSAhdJ
rT7uemSoBT+bqwmCMpCIAIRo6eGv6mNXStRTGne4ux60hbz9D7Q+ylUDQPRWSk1P
yZE93IQ30P4I9YdRFTlkAqw/2ezhNmI/LxKtzOaLogozrqQwlyeupSMQexzewMW3
cV+AwTNPEPkoDraTfKo1pR5LrMy2U61i37LxKRqu9P+czFh75nVuT7iZxJGXHdMV
sUr8Gs6d1T3h1UF6i1qrzPFhKV/HbsqocXuEFODL71IG0i4OLHK0hZOPpz370SIh
Sgw3Qq5HMEvDgczg6rwk8BDwrULWA/id2wgZODKotZBh2yq910C1Ku5DZk3NJjRL
1FsUkvJw1w3YzlQ8h1XcPp2XQbYYd166Z8+EDzY/Unv42iLPXNvWDNjZFkQ0cI/G
T6Wo8pSR9/CzcffZ9MJVY6W59ubybzYoRf1jrFisVm6poR32IlBq5Wdm2nj0WXrl
3WG/emfkHuj9lzlCVOz7RW7dgLltyxFKnFqgz/j7KUnAwH+z/rXdHx4Xhf9b7W6j
/5zTmiFxopBEV8UliMNhud0kLHy8v9kfGt9Fsk+VQU5kRSO3HqJ5+2FjelzBujsS
HqtL09dYeMZ7pjT3+r6k/91Yo5xi0fGTtE98QtfcXJlwVS7gXtXJLV3CYou8Heu1
q0e5MnBqyCXUKM/uqBKwBeAqY+ZucR4W3+82jWVg6szrSuTEQ4xkQi0gMEqoLsHl
MTELW1w3n4D6yO5YM/W6hCtV4BdqJNRyGA4+urrP2kLolv3sKjtvLEQ+HgSY4OVf
XbBL0fGhOnbAfBWKlMzbGNBNhJ8okMUviR7LW4/AT43k5dXBBK4m6Shr0Om6G1tM
xvZeeFq0038uyQNfX+X/MhjXrgtY060JvTXtPgY2NfbbCJ9FsO7UQic/Q1F50IOB
P5MkzDV3cGSktae2QnSWpTREIc42z2w0fJDS011DZ+Co3l5bWXQyZ2lN7jXX4jxY
zWBRlEy5u6DGFuxL8wu6mmJ/iY9CSt2NaKRze/WIo1vaMS1RVLbuV5LofhT+3oXC
99UHsT10QDRX9LKV6CAGqwckktIe6fLrqDQBUZJeVUP4CfNQVcRJ1PzAIuagqhHK
rDLqHkWe/LJamGq2dTQF93ZuTWv1SWyj4gqTjWKtKeo76W97CQLX8j3u75fgwXws
JX1jfcstjYC8ykpLFxSL5EHk6fjYdVAkvgua92CYN5U0x/AaueO/fdF5B3NMMxdU
ZrWUZG4vPyD8/at0zapQ5KPW/VhduM9zLqgfKludgc1SFoXIuYkwsWcjbcCs93SG
RWWs+F+BhPYxlYKvfCGLJXz80yeC40dg9d0NOe1e2m3wTApWrWmjpmNhKJp9CuWi
L81EHBWhqXAPTPRjUP+HlSvIgMVudC4Ket3xuIlFEVC4/JAPpE614w2bHIKspJSr
adP73PLB/hzgSLZVJp4eTRCc/XuUa1sH/I10qsY4dhSRbtYAgaSvYmag9EIkVV8R
taW26+0qf3W4hdQuqE2Y+IGqJEqpXuWWM9SoE9o7CrQ9dybhtkfrLfQPVcY5RHLp
ROiX64DtevmEd7SUvwDU9rzkOGDB/r+LcxafpiljjXzkPAdGPflPzc30aV+As9cX
BLrxFXpOiLcaRCs/34oMOd/W1iBUe4nTnVZKG1IWH0lL4Rr5QFTXIz6FTydcg8/P
gQuLeS3M68huYxy0d/vBAkBPPAzrn6oSa5oQp/ChL88gJa4z1bE9C5AWqIxbyPcx
ST5y/7yM9J0vRKRDEGEbcuXPdkNI0GAq2tb4zyNcJ3iQBK6Bxp4xshEakRdUMVSR
5B8oOFz1kUKPmclccuX5ZQbs3rgww8U/nXyfevDxl/vzRUQNfCq1no2hPRRJmCbY
MVC9iOMxMfHyRjAxYw+2q7oicebntyJHp8j2lF8INCwyadVNxua3l/wEGGW6J3rz
hpqZLzy8jSFu6aQJfPfHLpzQIr4D2/CCS3Iw+AuXL7j2/gvGliVRRIRzxYMtfShV
PBObemXn7Vpuo5BsBcg/GSu6uBgZ6JB0q5nM7QujkypbNUo2Ou8PWLhuLNpdLROt
TQ9jQUkO87RhDnq0w+NJQ3+tnZiAmjIQn9337cJnL5BnLwcVd/slrqoh7tzD/9cl
zrako7yMLQwZQgfKWluL6HJAV7Sf0cK0I79jl8n/Jd7A09L7YqFc3HSpyvE0xOXP
8aTY0ndKDlu3aVBhQkKgfWoer7UObAmRu4K2+g5+mafmzV+iantjJ4MrAvuWOWHC
+z0rjq0ToktsslAiE5eGhujRnFXe+RikkfKhxli1xYBLwn6kd7Q6cOuBk79AxqUA
un9s1BbBG3yWClHjrKZRq91AAWQaow4tDixULNAdRxXAjzdW+RPDPUe3BGCFGenF
c9wwYU0yAPmOsUWQjoHYqdbP+wjAVrAZOgiPLXBFx9NFJUy8SRziseGCSWchJmve
wD5AEseRj/BdxNmFifq159OoDQo7u+cHjNaowMdZ5JtpCyZD8TOZa1HghkShMVmR
QyS+GGzM6OMTpWWOR1cYZlEmLk75HcsCbQtch91QR2NmhHrBgu8cJeV3qMAYnhDd
cn9Ep2pb6//U0ZUByYNucKcG0UTzGlPpsKkQiR9m/NbJrFXdU3qHZGKBdYX9FpOI
2fQn5wv6o3GDXG5FIOY72df7dYzJWhE5JRK4zwB7jqR5DldaN+iJpb2CRtstcIXv
k88uxv0odmvnRUZBayGpJ2HqLZ3+K7KmpC2sp0NpGx+5mUT7RhEtbzf1p+FY1c9B
jUB3H7hVzj2t+v5gnoGHfKKKbJpbShoKf6yRSRGRNQhS5aM59Y+UElgXIZnLxvRr
CjFzgvHes5fXa7Dh/QqBdgx0SWoqTh+XepOVs5Y+GvQi7YsmyGrp0Q0jtfrbnGks
bMOIfev0+KMuRoD2HWvXafWtyfZZSGoSdGqZd9+Jp6kZM30HDbCG/VGW+AeGZ8mD
LoNTrQwE/Yj2CGjxLf10imALgbPVlwLN0IQA6tg1h0vMGB3dBvKtQ35EVfwLrKJu
dBALsZNEYNUD97MxWGoB+EShi3uxPT6OpBteU2vinOk8PNLZu4Fkt0Q6zDLcinTN
53wLMVHUsFG6yOUqzdVsgt+XTfhpp4aQmUg21qAVrfXUOXJ+4xrf33xpZ8a4gbBf
rzcL3/K8PtE78FEf9ofiT758iWf4lES5zrLf3gsk5/1de90kvPqkXlharLsoFVUE
Jkg/QkPB1VchR3npbtIKKT5KAbCfrZjLwc+57nzBjmbmqvw4vyz6O25DDPhAXg5P
3QLxqJT30C7c5pmaVHXTOeb5ylSWgO6Pef4gzNaNX48JNWJaiPZee1IR6282DxxV
3duR6X5Jd1ZvZ008lj7YYbRu+2LvAk9bkY2qKibyE9EOKaAcKI/rCx75yXEhGNSN
lhFyTszfGq5k0cfsSTuOXiLMKZcYKcNWbNVUAGoqjY1q58urBiEp0a3of/3j5Nn+
7y/L26w5zhHHDubAZjZeS+FCbMZO0I5m4ww8gjJCQuB6IrbBbgBvCouoAROjIPb7
2+2G14EyRpyh5/IZpeaya0DOkgMCEltRUZuV2OTAfSNA+EXJ2GpNcwLKEE/MagH6
76hFRld1DYOthBC3Fvi/O0IHxS4yBZVd4e1e9CXlVkyIoDm9fgJleXiDVmbrsFzf
05lTujv2Er1rF3zpAi1FGhl3g+PojjyFeP3XBPVrsCEBcFnkShdetHhfT++onI6j
nOrT5BWpHE3tHnkq2uhJqB1MDTMNJgTx60Aob6VhGXMv88TOkLybRErxYvRLTReD
SfMAcjOxxNXq+PlbLA6yY/A+rbcFJmsw7UBHaXRMUH2DfOYf8Ca8hmeXpKYfuiRA
4NoPKD1Q0w0r1Wg9DnTNFAuBNuNdPJAaujZ7ZV7yCHUCO8OQAGmEC2d4kuWd0EwD
+cc1HtU7EhsWVlUCR7PHWUGkW0U0FEOBY/A6Oe2uBbotiaxFvgqqhJHXIOPzrTzA
J+gUbNoTyVaNEXiVMBZGS0Mv7BWvol5lIZeNleiZRKmPdvAe/a6WG0ixZJRHfp+9
wDltHH3IuJQwqI1DiRldV83OErslETw0k1cynCLgCpUVxeC8dOst969Q/koZceKy
iBaatKXVkyEvvA5snORGOZDPJd4lGX0l6qjLD0UJd/tsk4QS0XUt/qYcmN8XNXSz
OevRj+6XviJCftDZWeH5mb3lD8JD4H89cXwjojNjH5YL6dTN83vE+4+9ce9p9qsf
NDJ4KvGp0wxMImOwcCwsa28ZMeGmFg3bk3DKeX+5zVt2sD/UzJ4No+UraeteM6Jy
pUV1pQBxnddJgBvIGNAldOL8+rBmMCyVT4pG4sQJdExJSkGAYBcv2uJAXT7oGMY9
AOrc9e7SogYYjfnBOIox2cB7UR1VP1fJJ+9C0dV/S3aNDorImLc/T7vTogkMb+1+
lctIOBrsP3bFGeUEFPlyoZZCKY/STrEgqPzDYHZHfUJqCh3KF6LMa5Etnm+KO7Rh
04rn4N1w6tL4OxdyE0oaCQ5ta7hjIMGEcsSSb4+UgoRMpZx4Mo6h/kWhw1FVsM9W
SkDhSrXl7XypblyYU8SO/Dh4jc7TABAFH1JEryI6I+eUZHtUxAcF85ZX72vsjclM
pBe/zMHToLIGleB/V59BET2inotTXsmKdn6Tvh5cS3h5VQ6bclNQQxZaN4tLF5sV
wUhdBavHMSOB4KfYbvX5VsSzFCrd1aI2utqinB22Q2lw3LBwUJvJ0XFfFdWgNDh1
9+jk4305G4sCIrI+O6IpsCcXccCAbVoReIUs8CIEZGHA7bxqbLN4lkY2V7MZq6rw
pehXGtZGtfV1ACtePUZ3iw12mh8nQG6BexrwHmxP/T83DcxV9p4EyPOA+KD+m6ka
TrkP3vrdG9suA2BleX4CstwsVxYpBd7J4eHT9Q9cyZveLP58rJ3ll1Dc1msFD9LX
nC6SxysjUUBLP3uyNcM8QO5cZN9M4kVNUkI99/z5mae7JSM0zewZJkin3hpni4aZ
U5lCHcNCkdLx8AP/lSYrmlyvQsv0ecmlgNIlau+0+52KEF31AAvnCJPvzP5LSe5I
prkjwn4NAss/6yZPi9dRyJRm2ctjMj393L5yS8U/u8mvgxzzbLmzO6IB/B/wqXAc
cIuLn06tcp4QjWFNZmGNK1GnT2uIAGt90xvETlZEpu0t9Dt+BEQLWJO21h4xZbry
o4H8gLV2xDh9P6HJg1qeHBf/FLky7ni90zukCEshKhiAjcudw75sdfWKojGQBNwv
phLrKrLuJ3knvj9VKOxR2RvBYEKyHPrwmkrLuTk4mJOHgrAYe6RfcLTCfn7XO8+s
5fSv3l5XYgecYUmoEoNi1ugO1zYFh96x7nDr7o4dRkCgTm3ftwfgZtEuNnKqNy5T
G+oqppDh70WgPpgNZ+ARVMxQvjygFN/QBPug88CdrBOnOB0O+k9v5F6JRJvsFAhN
w5iFvgrAIOEoHK2R4cXna0vbq9kaCCk4P5DbGlZ60SR/I6C3EXihMe+OYOrnZCre
1F0w0bozeV32dMBNw9La0EHxeXEWPT0mJ3UEar+GaMfWOAQIYv+kivlbfsVXaU7f
+ZtaASjXbsX2ygjwSe1JgBGkl51bMKRwFEjtv6hXncalav2MjHcUn1GFVn1ynj6U
XETxW2XEa24QRPkLjmselqCzjmLlV3/GE6maEhqaTuXWStZvj4lYbv99PD21gpX8
Daybv21EqpBWVPNxpCFuAQkqMlZ0x0hxb5K0tkn0D2xK96RusaODnrKFzeigf+E3
/6MpKdNzB38zSeoR41NFQu0WuheWFym9+gOAzSfLKDvs0eDa1wg6/vsNoPEay06W
JXQ5FfK8ZgCiIQCigPyQFWwbX9U0Be4AtMC0o35DSNrrNOGv1GvXmHhTpKPZQu4G
Xhq+x2vEPxxPDvwk3gdNMUt2O0yzTKQEQHDxcd6Oc3so3PwCYOtCUpYOvSdTJeHk
3TUq5unN4USAosxRyRLrbyj2RSZGA1jnpySROVzHpi6vW7pFkOsBvB92Xv1wJ2/k
ym1mq2aOu/UFuNLiNEV7yQA1q7KqREzlT4LJMLndaJmBRhCQN+AWpOIcTFxoYMt3
WOu9YL6eSBwXwKMmcJ8yRIvFI5beyz+i9AdL1W5mUEx2P/4fn/lS95YPnLksEx0l
tqsegN79MaCw88Su9AWG0Pa/oxX+xsfmuyr+soJS4dRfHCcJRmvp2Fm4V0Mjta+C
J9sCatSI7kKakptgp+LJmWi0lF8YuOG/4XKYpFKcKGE8xiW0QTjBLrPmlj+fVaYj
rNcVnL7hFJmAiS4zTtDmxxQ4ail+xXPdErpn5O6w36Z75DMklRdgURJ3FFpA/9GM
trqt3/AhN0pWHihHK5xxkpw3MJiLtUiSVOLYLqld42TVxwFJlDimJrb4YSaOQzaM
oQbxrHGuz8CqqiO1JVlc0qzwLb2Bywj7y0A1L5K3kXiqkJJw9nNeq0FH+tsH+mL1
3ADuGEZIphKIZbwAu+m+1rxcq94qsijVWFrUtkJA3lFi30Q9Wlf7pV6SkOV8TkxS
hxhzt90KLJbsUgp9Oxp9NM4sAveQ5FqROzKjN+q19GDUAw6PeY6k9V1QZ7Lpdojh
fcuhR6o7uDhBXGJZFuoUyGUXFitAvkpsSr7zQMhc3rYwj1chDzJvLzaDxul7VkCB
ScjrCO2RWGvTImqGLHEhkZFBA60fM3KlaFu3JDvv5n8M7/cmpPeH4NooDrDgXYa+
Fq5nBrY0HY+WRLBBBhXQojxl5KdwuG/9wNlbwqluhHZPLjo1ZZnT4xxuyvfDzOM6
V1kmrn9lWdqjYdChjctd0i6Rdv+Unl/ravU6z4iPjj4tjpadX6wZTLadr6M77sED
1TSK4b7eYA5unr+PHX+bkGXkAC6+A9G8bBU7+MhPA75b1CbO3axUFEuzxmi+iSMC
1pp6j9Obscl2iKG0egMw8RnipJswmVZHxUCloUKtnHYvEmF9Xt6a2mkR2AjdTW4m
JW+da4a6VQBGqd/7F2LCP1HTaEikQVYkWGTl9A7k+C4HTWsIse2uEwWrRDsUI7Vq
Au5qptW4LFQV7HCYzz8x+WIOhkiDayg0YK0J9XC/9VCHrc8Hh74f9T+/SmCbKSD3
f8HJJiOEsU365CjiDePBjZsAeASWcYKpyou+/WhyDGr14OkLU+kQtXSh0M7ZTZi0
nv0ozBmn//VTmQgFZX9/SXrF8voiKVnxs6LHEWUdgPB/9KrQQQWU5LpAhbjIXYG0
i6e02eeBfmZtTfr1gJTrBlh2msk7r5gOT8vE5mD87rL4GTxDH+kVUnVSE1SzYiVC
bPm7mR/0X8p3cJLMhfg2OLzUR9EXXkb3Bv+DMC8ET5qeaOnw09a13bybCYKsjN89
PVhBIk/HWSCF4U28zKeshYAbqzJ7lbuZE06YPn3m6Bmbq04hJpDsfer00sCKBIx8
v13LDhuCA272ayvTyu2YGt4yH3TijJn5lEmLK7dg11PXstFIDcLitermudU0MPu0
ZWdtOcy/YlMmyRe6D4fCLRMADe+B2i2BDXnv1JKNcPcM+VCOWZEADTIsweeVLBtT
hvF7JPX5B4JvOzUowQ82LWmaZKofEfE5EExkMZNSJ8Gc+tIMQiF68U8E3KbKDdkH
tHz9MFTfwAv6X75jqezCowZJTDaKwfZPuLFI+ZIzM+3M2coQzdynuOQQ5jorp7+u
g5fovuXhzG5Jgeynu0NgHfdf+qA58uJTDAXTgOYYm/VEMsvaaAtlKa05A+21TMW3
netWBZlpvZ74aIytHVXB0VALWhIGi6T9mB8XAgwhNSW9ze/2RXLmssEFmA+zY5IU
xa3zEtR0s0/sduyjCPOoDUBgH70vp4nIhs/AAUmemBKr7/VQywUFgdJJZxFr9tmG
Upb24GQREkm+JDEaT55yLxukumT46bu+fQ0Ze1o6iaSDY8t4qI+x4UwI0V5ODFLw
4aHTuDTU+KxfY00edDSKXJyGFhyW9H4ApVjKQFfaprNNQrgK4shtxTFzWp3EQI8o
rsfLj6dKWfGw95/pxdQW5F07YbU2q8McxRn1zi6nQqMtPtuM+uWkH3mbKz60oeI3
6KP0dJhE2FRs+i+AgszC5+XdINRam4pPNidBzSCVm5u/W9/E+P9BZ0pgEnvjwbMl
IrXjL53B59kc7Gem6qskQLCepb1bIq18P4bnijGOnWhcaeG90U+qV0BxekLVAngL
g43P2gL32qMcW+SyxWOrgE8fGHbUdd8tQDMSsbWDcdLPqyhhx5WOjPqqDsvalhbx
Q0rGfTFUCojCUmywu8NICYWHCfANY7qGVSicJo5Hgwc8w7B2ifd8oGZCCCV3/Inu
1yqIPGwQSWKO5ri3yh0OjHu2hqOgWiRpkLN4w6TYTAKuSEcUcdjned+92qaf275+
8W1G6x6spf8f9/E4TFdfHoGErUAfDzr3jqto/7BFks5/kNlir/sS9EooJiGZ5qvI
JUOaLMME04twGHqVbfnhNrCjHlX+GiWs7kDk3oG69qn4u5+UWQIpdt3dtf4aEtxu
i8Y+wuWRr3QjSJQdyruYqwug1xnXqB7EmYY1aOj6hU03a3Q5iXb5WyQIj8UurLJl
ISrhNuLjn4Beu+feA0lyTP+Dvenp2nlrfVLXd5j+43LVL4Jn11I9exCvXf1ZKui8
5iqL6RLmh3KeuaV9uJhVu4fOAOMfxRyx1Q2WgKlR2hzxg0ukQiqpdfIT4ZUwzUJn
7R6uqqQGxlwGkcPS6IKOOIAcU2qvQDZRC2DHz/1XaApEp0dTD7Iwd0waCjYypidm
A9kF7q1uEaah0deih7LH5cLnWnHusHNLGwuQNVS/eqAZ/va0zDB4gSVVa2lWkuEY
PBO23u0mw9DeAf8bRS/skmmB0gPVpOFfUOH6APERkyXIrnzPU12Id91I4Gi7OWge
gXNOMvKJK+8YLJNh4foq2MZNWW/rr0e8lSLi1vxDwqMZzsvKSOYmkktJBBB8CKH6
W/rxfjk4nWWgYKzfxi32hc0UZuPGlf/9+uo8G5lC0uOiodoT0uwUnHgCEI98q2Ja
1uHZn8Wmszp1fdU2J+svz2050EZWKQWntZKfxXntMLpZhZXbRdAV/ohWDWjoA8N1
pX1DIEGHQ0QsB0emkumEkN4b3jJGgjhBMEqFOqFvOo1cfGwDOBiHRVXNPyTyvxOH
uFGiwwgiXTpcMW/edCnVIEuRam1NjK/5SA4j8J2qo6PYL/Du5ltZhjLWfqYfxR1H
nqvn9L4a75C0q+w0vUbOp8Ri8k+0IjvoPpiuZOjBIvC08a6baed+rtPSru1UAwgn
mfJOJ5W5gf8uPDKVsvW2KQGc8ujeoaUQIRF3G3C9FIVm3uUcveXTxPB8YhMtuR8A
2eBBwpm6fd30vmRPXaytXcDvTyWdUcMBtP4KQdhwwcWz86HZeDGB0WdMFKB4Yb2B
KER75GJXlGvmAtDbAW+UHWUtPfq34O1ddEy4+sSlfgP+UnNMAlpP2ggngPk6MZsc
ZRbl7+B+IE70okkUindjPMEja/ehFU1105OdbmtDooSaAEptgxi34pdWVeat2CQW
VejZdyo/MpnQZmRWU1lz4rvn1/tiMpXMyCn2Lk5g0WGmOHxgiUbbb8iPBf+zTOy4
qgp6S1mlzbBXwSVMtEuixPU1WA5tiWPsdnwelaJUMkIUWwNfhAyTiCC+N5ZaoELK
whV9SEHVLY6oqMVg0bMQkwergp0r3mctdClrVfVJXZreom/ACL5JXYwDuUouKonZ
vtY3duza7CZuiMGZOeozzV3sIOnf2JKm0xgFklitqm+d3CUwjJP9KK3AX2CDnsil
1oRLpB+bV1WIIGAnEDjBvdiOAlcmO43DM/2QL7+D/r9CcGlK4IBo5tSH1xUpzXoJ
n7mJt7zV/QQercO3wAV2mPky2YDGg+OOkm9/yr2cTTrh37Rl+N8xB/n5HIbUeCzJ
etTxcL6nAH6XVrCIusiuqqiAg6XzOJCeqw6WF0kpdEV4pK4WXDjE4pnZok9Co3f6
RishkFtTF6GrxXYZsbEAZB9lQjcCs7GYXji/ymMl49OdiLCVYWLsHtXBgpbFDq2b
7s7B28XLbcf2ozhWARaLsIRkew7hEbHb4WAPVnJjHBQMPwECGhe7GTvUy8n+ssHf
I5Wd4Deij16BsmZfhRzEusFHAUBMrZcf1i0o6qO0ls4pN+juGv3nGHO1HzwOfa5K
65WnUQ4PdLHu0wPCCj/QzJiqqxHRrU3YgP3rj3O3J9n+Pj7qRtzTeJk+1VwOXCGt
2wGkiy+RGVPI18eKo1+Guj1vBB8s/FpP+meZrHssUYnEqZPXgYT9znH/XjYcuTgg
BPRBA3hAP/mRjhdU5ZPP4aUIZfvlKhSSGKayo4xCghssK7Eaw+nohshYYhz69ea8
Fb1JccHKmYdGrSKYOhf9dXAdzZXGWbECVZ5XW7JP+CJTaaR5u6wxD1q9MBF6s026
dS6A0dCjr2EQo53Q4n1WCcBwoEBZb/3y37ncdXh2lpBJN4oB7Cx695MLfrsEIagp
jG2JhNbkqHmbd+qi7AbVeKyxH3CGY8n6MkqOzTHum8psiaKCh45T8uPBUVv1HzWf
qZa+HoU1rJq4NRBEnUqn+RYD/o7R6/OYW8CuANAE5jb7f3JWL0T/shMnEuvJeLk3
8pvLh7L9dTZbdeZrdTIttpX7u5+nx8BTIQXHhcEPsJ+nC6AVThWtZMuBHNVEU6Je
a8CGOCEhFvb/gjqOu2eD9V7xIbVlAUmCsYYxMMypifE+Xi8IWevfkngT9PnSfDdq
ioWE2tYRA0uLdmP6UeRxP93TKFyuZ1i0TkTj40DB2awNEufu1VZ1+OeWCMTU6M9C
28z6E5g7d09BApaRL8NRqXPwTb9sheZRIYCK03CbXfYq+YEO5qkowE1Rddtk3uQD
e8oTshl67gQEPmzFtSpU0mNWcQ3BzhqZDDhHwscVuXXen4KCwJ1H8jQWxFNAEjF1
eANA+2XEAQdQti/NVm9U4XkKBPGv4zoCH5MmR1YqLuDcQuqktgAgsEEyyVQCsljf
jafWdRHYUR5QIdorWCOYOSOB+YI1k8JhPHtHRMa8WkVDN3QCEIwdxdoKsFM08Bn5
BwaXgL59XQnZeKetpPRTiql/+5BtOfY6nzcdcDjCGGrcMVVr2lt3X7/cZJf77dZ/
4SAEOez9ABJ8pZLNTBp8SVoKSM2BkLhr8gkK+kPaF11Fz4TekN0HM+EKiZdeMdoQ
+Vh0ZNNi7CyqkQ+stIL7ne7PoEbsqmDvOY2s445gOVuoW5/1nxmmjcqEVBtMo/md
gh2i4lEEjk1QcCTanB0IHlm9nfQC5k5ds7iWb19c+qKD2tnXiSuzv4FDhqo41FW0
xeVeCNanpPZpiy7Fbe9NkamLfLjHLjV3w6MP6vXICXUMJz/rYWlw/WCxrQIfAp/x
P3mW7gm+4H6Py4xrmUg/MGFRCbz/y74DoDH1moWw8ysS5nYNll59g89nLcyTw7rh
Q2LkHdduZJOJ5mBTY/XQEd/YZxoUP1FOE3VP7nkUu1YgeXKKtdBdtD+3ecJRyUVZ
XUaOiwanwXzZGtAL96p7Akq3U2GJxxvStlMUKod6MJ+UovSzTtzBO27tM9SlXQWe
p2ATKQS7MQdZuB+uhkwu+JMzc0MbuRaJGLhXztZtSMK/LM1+JXR2aYqSSpyVfwDW
3UZM+0ZIHdHBQ8y+o7XKN5GWwp448woHqRPxbFOuTwxPwPp/tiY9CqcBsw20FXEW
aXyLJe5r9aO8ioGHhS/QpfzMzo0RXqGBwYZox6Jiu/9WMlpagG6RRGr8RuzXlEoN
qMwVXh0o+W9d1MkrMa7b1KyebVIcH6wHKrrCVechqQNp4cG4tz3p8TXiyQrVwT17
ZZuYJZ6MRFIMEsLi7t6VoaLAlYbHNqtFNrcsWMcLf6Kmr0ogKK0DVm4CvjSIg79P
UgMHITUdjpf41W0iIWyA7OoMw0S7yCGQHcuy26tPANvY/bSIw6EaRHBaYkfu9JEw
D77jLCWKgYDBDc4KMzOp1ZnHy+dUAAR7QdaKbCnXfpFMhW3JJziE0Zv1d4kKvoci
+mGLJS8gRdARiqoaKrfYc5LazQp0yoXWRVbLbfIMJyCqiOn30Gy/B4d81w0210MQ
MWXekgQ92KSkhOVqSz0fQSHo9vvDTGCsHyF/uN3BkffUvppHMV7K+H8UHKfebr4M
27u0hCkQS/9hNydgRgmt7H65bH84v4vV54vbhPTKKZ0yY7xDlgbrLXYCi0TyNGrN
YkkhN3Pwyg2Kh+Bxgb7HKsBI7a/BJV6h0MnofKCoLvNiThJ7josyFD/NNvlL6eXy
07pRxFQu0xYQKXFASm3VNJIYXvPckyQwYyXfZsmquEEUDeeOco+3Ern9Uwg0h7uy
hVJWBBnPnGQDTNEwZrZOe7sHKnmkRS59tMuIZ7GGKrZfNOfviWL+YzEuLIVgllox
e/5xkqrd4wQxHyv4OYrWeONIQ7dVknFfMAz2Ojwe3kKCfqUzZ6q2Ysosq7VHgTVX
N4yH29mNUXYoSJQtColFBArq0oWPyjdwNaV0krB6gcDMMCRRjJpb6rInAksZ+Xo7
DqIfBnCOXeqRM3STvIW2WhPu0FDCmDCyr0N4dmiq6tmSRpo36wTBsI1ajiw62qaT
XbAChtilbLuP2EusgGjXYCJJRe9SU7BohkWDm4ykuCB4fBri23v5tvW4HoigFGOv
yVxEdZUCH4qxotMJi8SOyOIEMHYNi7uIaBkMkD8VzgoIYYLHOJTCw97C1GpmrsRF
wIG8MvEw2iW/jFA37GGIH4hIeDw+MgcCAlSjmQ7EEYZDGWCjbG7ICdHIwC7RJaUo
kRNDYN4cfbTXj57xRvq/E8H4D1LKuxdJM7bO7BabU/d0Cm32UXs5mua5Ul87IHFO
2i6qre119mPSYR0xz2Jdztimdh5AqD0E7amT1aSafhstU2PtM/Spl0JVks+BC9F7
yI7o7uDpgkfFXDe8tioObVpcMIMIK/ZO9LoTo2FmQBNyzQY5FckWsd1AmfCsXnbu
BBgUSsv9yJHKw3IsygJTdqv3IGGi3WuTdLmA2n82aStPKxpt3AumqPFp523+QMk7
6BaYg/hLHJ1ncfb/BxqLL/S2ZwD4BT+qOk6IxmfiGoK2j3/nb+AB6U6/x2fg4xdq
OusgleQvFLvIPCgBZno2913SdEvR3Tjq95FJc1mQ0HAXRKWDlKyd18gAiPm4fD+R
3wg79qseUfio4V/4jwDncBnrNxokTuwdtsIXDYtOJkncURs2CM1V4BWwrnGgaed6
EI3UQThuYncAHE3gJ+XN+yxFtVtirUHS0xX+QiUNPDb7s/Dsrwm8+vCn9awDaCqN
YPSK33qlNqFqSEp4B4+YaR9n37bUqo1xusmsO6qLI6dw0QL9J9E069IAq64bwtlu
89rMNDf3AKDzjDMpsvzyngwbkOOr/KJ7q16wRl12U2lxxSkPs5kbHOKF59uZerr2
/fCeQpL3/bR/chiYw9wxTMfU38RWZ1C5mVvcHiVPaO3M9EIJOc/Z6CU8eLbIcZ/5
E+z6VYFL8IldNvk4wmcNzID/tzeMHCQQNPyJaII/3asTc62+15fEWxOgaoaB2x00
Rf2yq+630CsMKgChFxzEbUF7/MbpgwVtSObjozpueGnVNba7M9XqKQQa0Bw7QBHR
k5iLd6rdiv2wEdO2VxIlest8bqh67m9eFJCQIGdVUH8Qn9tFCtc3MeDCBSfdPbFP
m3cFcz0SPwz8PrBVqP6UsV2wOwMU//oOGs26ZnOx+VedDlgyu9zPHxOtBiTOM675
eHxPavcc6yXqOOmZTdutXM8NQZ8acwd8FBOM/uQlSjxT7DIeGhUj0DF2zm07HFEc
TRtakFBBjVAtJ+e+gWxwDYW5YsY8RCjdoHR11bgYCVje0DnOBePT42IsAatuAOxN
yQp3dlQolPKGIBKRGawcu63lNmmkDM8fdoDv8JEAmoITheWgUkpigIGO4WEuXqOH
9Cu+dDYrWCl9qdaONon7eoz1ixsm60wSiuW2vr3SWXMTraaLykc+s0gt5CGjF6QZ
+xwbyxGWRH1dY/KCr4+TdUHHgXnwOkMAZVeN5Oav+ER/tsnE6lJwAdUPuBO6bswN
RDHQhFlJoenYaVWf05EvYK64BgjO7A6ulA22DO6G7O70YFJZSBvnFSrG3YywAngz
ayEzb8vkE03cqW09BJgLdM0Ui6emyLNm9mYCiFnlz4PUT1/yMeLGLxUfwF1fKoCv
rL9QzxyWISBibZTK6BeMLNCq/3xmsXY5f2rny2RGV2PEFqiTpmf7BtIjF8o9vY8w
bWQd8nElKjqQeBpkzqgSvDYwq2Ny0l5E/zcLjPuIA8Nui2M3YK7gUqmPdnun6ybw
rhcgz/cPxz2DIHofjmcvevNOKLnrQ2luGVUzBhnHnBbGmbFDJpVlG/OZ25fsv9mF
7H++Tb2VHRJme2A/xP/RU28FnstV4vOAmxQZFP+sBWR/ozA+eML6NcCm2lto4mNm
NIAz3yJnPWwYHZazdzg2tTpHShhLhshnmBFNnww3gG4FHZo75ul4/w6bMc1LbJXg
i0RvyQq/wC13pusS+CNnzvDYUE1tlq0Rq0pdsjkjGoz33Tdl+wpN9h1Ky4v1KiDa
omNhxprNdlzYN64eZeqSfC0ImLHxROkxM0I4pHuPoB5ZaJelHzGnef3X8LAsQx4a
2dAWNGZTsuUROEMDMYZqm+z/wpNtVHgqfIckhuW4kqdvRsvaFSB6SNy5fxBbVExT
b0HqSN8r0OkDhfW8zbROzB2ZQRkR2JntzQsLoBxw+jWnQxemnqm5kiUUSR9KwoTq
XXVPueXVXVYfysP0lHX/nXNA08eJ+vQN1HM4No12miVUVcWWGU7TvWpSgYnZmyxU
nDUU1upXJ/pBMWtZO8x3ZedzzNrFWZ7QdNWa+vkhU4Xz998TyCPAOzz8209um8a6
A9AsbHi0KTxnO5CD0sjj4pLYgW5TWrvpZGZ/L8/9qbI5QATjfKAcKQbgUB542PF+
EDfO4fW+S46tvM2FtLnL7GKsrxm+uRcBSYZEvVxBBsXtf8nOLDRjorEhtGYrNc8H
jrHGjnf6qkWlb9xsVjJpqvli//rP3eLcHStIpU+oxtCpUe8cxdYgCJCST8O9BMhs
D7ZDlXCGt15ikisrZGy+2UiSkMKLD4R/7qg7xLX6wgEVSd54VvkYrY2uulM6cCbg
ZV+0RpILHrwpnyxYZGSsdfha3szz6vQ46vrH78tEbr+pUpTnqCWjbEdXHZLphCKr
3eJxQbF/kiZsdiR4hBRkjb5tqBbfp1bZNWzU/h2brUCcUeQLMwq1lE43bvdEdifI
slFlbnwPivRvoQR97MZPPTVHlOEh0LJviIQb1J86LO7kq74d2000sgwEID1X1nAR
jeRnIefigZp4+G1IrFAq3CEilJobG4YkhWbpa7F7EheJpt+B+HFMkCxXDEsOd5w6
uOcRLqbCQ+5EowCWIU62l68Tg6edRhUf7CpuhoKB2PX01cpBu1nAeCg5PWKJP3aW
0UXMyo4/Te6tlvo4ick17yw+IrjD9SUsem2Zql1nkDVI67Ic1HRAmQjtck2zPcyg
IYGGdOed/OWcEzcCLbF9flHKibqa0vHQKkN/o9/jYJUcbrYU80TeBhr62P65fUGU
UUiqAVVjKaFyMybXBDvhyziwWBfunB2ouu/WVzoPsIGHNuFVytpJ9Tu4ksONVEeN
fJFENZvh9GPwlbgUZZOKKqv+u/I6y9Qt3fK9Lgp5LYIYrzrO6CxxoF5LcR3hcxK+
LvaLWAcglMsVow9ozQHjQNcTOCC21ju1ZhrhaAqIq2DQPhpx8UooaEOKVmuzzY/O
jBbovck0UG8vmhgTxkfQE4wmVw/scEXXQNsj/fOYy6Pm2yfrfKa3KNahasCTYLYP
LUgJ2EV/Q7EpNuOmDFu70MosnqE340YwXAyX+La8tl8sW6kiwXhrVpYH2bBrN1SC
Qm4eSdXsAf/aH1KY5sAnAhCI5DVubk8WdIxaiqdwI/tayv3g8o4vvZISjRErr5bf
pWdmkTPbmRKlGNYz7/qT3fJ9/Cw3jIsMuTuvYQqXiWu28RdJ+KalGAeeJyn0X7Re
jYGI24RmFKlZKS1FMa+CwX3U0A9nrrgPhMFA0BFaUeoFlxqC4bAEhY1QvN75HX5T
I35ERdUQfJB/nRxPcq7J4jZqdkfpHtZSlaGE7Qp+n8ScurRXUMwsU1JHXmuPwLXn
CdbJP82ZPUoG2WN/noMGNmvaTdYaMu3Gc5VMucofJ1ANOzep7cbXJnglwl7Oo9JH
7GlcolKqHaU5gfta8Rm0N8z/O7RXgfZkvAjiQJs1bW4SZ4qcoV21mB02aWojBKwl
gC9Puta0JQONC3j5u3PwucwcWNwGs568MU8es2qd6P9yRt0mBklOR+k1rPoUt1CQ
SIbo+NEGdA+FBwEtiv8KVF4ElwPvo0B091HA34EolMGQAjm8C3F0Vg7ufSAJpQHX
8d7mdim69dKTOQc9X6k/tVuSRWvnj+01ny//Sl6AP3Hh//zNev1VF11eKjiYIHOO
XoSAWexettv54j/ovGEEpsTFVRu3AHqGZASyatr/2HxYsFc8InjvIATnIW998iDj
2Y/GfleVviZuTyw2aDRV42Q+P48AOHE5l0HGYazmO1+vUVNvbShQxvg6FT9n8fNz
U36/fe57MEj4G+X4NPiHoNPVaNZyMw3umL3Wd2ilnInySdPdmihQwNiYWe+5r3Li
KkWjveBZ4+6LWlS+aJ2JQr0fRQV/g1fvz1FvshqznIqWM0H0eYW0E2fo8UI6V/UQ
p2QjhkLplOVwLxtful7zV/YFKcaiN9BLt7tyyjQUt/uOyvNnBGgFqF8C2sYQ4Y/G
0/zOzX5q66ME0MbK+rcSN2BVNG2mcwj2qm76ZkAMe0J7e7ElCfVV9grirzEOwYS6
n3aZnYHsaZN50Evxx/UifSdXQEP8iU8r6JEEj3nzQp6ZuV4tS7c+wXkbBCKrj5I2
tP84CSttu03BfSPBPnyZYy5EKc7a2vpMhKz/C7f4XaQM0QuVaxu/0lje0F3E/w4b
a3U2mu+msHWi35WyxSOHhV5noouo3ZqvtU4R4ZqJC+daDKsF/uHvfD54ZRI+n4zD
/n8iCqu/M0gDtLMDDdq5xUxGZhypK2QdtiHm8iCPV6nhM66DKEa1i7+WwFr6vAq/
ro5c+XVME9HW2oFzhgmRcPoVfa/pPpNzmZh8nIijVG52qpj41s3g7udNRXjP0QoP
eiqMQAz7emjrTW0JMSbvRLgUwq+Kw/Sz9tsXXLalyHpXSNpZ8Rk9S9eyaSGp7tAP
WFLmRM7B1WOb6mEWXshvpdlGEXmI/Ekr5I15vseVvMVCCKJjOguPQFvTXTwFv0i2
budP5hcWZNtVclZKwJYNfCwRzQiXYPWICmp04w5fBUCgDftYfXzMDEGWXWr4I/ds
A+4ymNOBhju4Y5VNNSmz5UPmH1lqkzosbQU7GGrGX75b5NhwLZv+u/q3952P50+k
lqnTc/uxLiLTJ8yPDChRlXIvcAlxUnohFMiDHH+X9Zsf5x1Q5In5EVpjGcjdiO1c
oVTZdiVbXwbAuQsaSWHz6jn0r5ZJit7U9HtWSG+WwmSH1T1hYkdm0a9H4nZQf5lg
2Wzaw/rxlVwLqPqrvMEJfwQfJ7zM/DQk0c7h6qC8yNci9ENnjtmUH56ws8KCoG7z
YaKb8pHv6YG0OMngUw3DY2/7/9FLnB0nfgQlKVbB+sLC2xr+tZOemXCh1exjcGNY
xbzUEYWqgj23so3NBSsLxNTUF8C5S6XGTNuEQZd1ECi3DTG5zCSM+eoMQcQoJFof
q/hD9As2JB+96wEXV6JBSyq131RYb1onVhzrbZGT7b3lLc6bywc97wqVB9rWu+C5
aEDrWNgFIrkA0o2jum1+HfzQIHuITVyEjrHZwRts7PbvbmmZSp8eCVMlh1XWAO1h
tfIeRhKb4iBalpHZhtNFQDbkhUH8gwQXWzWwvE0OgMG+8AiZhtCA01gr5QlCtUCl
iABhycfKE1j2YQpu+KHr08AxeoyYYIHXjGKXHOS3dl1R2QIdRLdqIkAoJjJ5RdD/
Z6rXd0re4+lIBiTXyCu+Y7BWgkJYr7LcypPrpYviyKgGIQRzrn4gJw1Obdugfcgn
HbjzgtmWvemLVch+FS/eIZDP0J0jSpuLSiZVa5TXah8LKkby/nHFX8y5HOlXEvFW
cD6xKyi7zZwyNI9BI8s1CvSuQ4NaCqGxiWycFCJpRkzTHymYA6xQXe3K039Uqzi+
a/BSzd7VNkPBMp/4EbVaBn/+QUOEdvuvbU55bxrc/NTtKnv5xiFjlLP4pRQRgk6f
Qb0DPA00W57ZHQxROhe3OAKuxkstJskVc95yJtSL1gjKZX0QpZnuoAhzJRX+B5Id
7zw0rZBILOvn5znSUQIsffgje9xvvYM0lAJWmwAwnn3dodRYjclHB/VmU87hkofr
gFLcAyPiLDpP7yma5nmAwTmhOQXh/F1N99kWFTiotnhrw3XVihMHKDYTFjGR4aQD
hYxhglCDDQTuiYtde73ITmeM6SAjgQMphqEaKYl4T8LIO6rUrXiVk+oq3qRWfPES
CrkPGNEe1/0JwIFjlNsCmBR3lhOvBH0w0+B3cegHGSTTZVkViQS7/Y4ZoeQENQo+
r3CRVrDTzminRY7nRDwHt00SZm1c2hOpRiWxFUGTOwBxtiJ62WufE5hwV4D//+tU
/Xq9qFbs3ZLCNnVZWOT7cRNtsUauhHJOa170WSF94ApRkD425ArySrsgrVQj8LFr
QIVD5Ri/NEN6C2fjwTYOwSNdn/kwFWgUKUP753hub4fx8Wn4OYp6whmBsvcpV5lG
40KIh0wYdlz1WGQUV2MqqchWon5GRgJ9fzg7cWzEys7DANjbGqOV5EIu4LOKl7nC
5UWeU2tVZ5CTzK+SUQMowjS2r5V7q9FyNW3skLcT5iNlDLaFA9Tz++sXyYINIC6D
3LEKO12zckFWh/J1M3HoqCe7MVzjosxmQZ2fLks3xOmYA+qa+oQpjK3MwYhxsO95
Rfkrj1q+ZtFXej7GiX3tyM2YStfWcxzn7rpBK+SOQT+8IXnpfZ1tSovHcfild08N
mlHXs7sVtUqxAJHbkAyfDSyaQ9GcUpcsbDC500fASMjgSYU+wFWYhW0PVUnfqNAy
HeqHhSiNzXuxHN07zxyZEGP8PWprLgyPYWu3fr+TOkISQHPD5OI9NQBt0+lJuwLz
z5hawQ+wxD8sliKZKMfI5d9w9AR8ML8axcRrPD7SgsHriCUnY5y7jXlQ2Udw+llx
b86HZDh8JRHES7pnRZ0c+M3x88CjD0IkqmqW3pEOfFCcj6hI9IY6ZO93RnY/r/WF
TveKUIpnFd2xzQTUawIUUHP/yPI9bSEdks6CWh08vPt5kM5Y5Qjtl2hVAMBUUc5a
PlT/aXbWbbzvoA6JmciaubcD3z/C8/HJ6qImXBaoFmdy9gXo9Rdgq8z/DeLyBB6T
vynkpk6+RENaSpY6KcfqHLG94tTlWZdlL4htYTJoIxiwc71EhxKoFTr7IhQ171+L
B81Fh6fx7sCCjPeb3IXhqKd7DP5UXJh4eXCx6LmnJNuw+JQjVAAYWjE2UsMs5PX7
AgY4haShosbN3XPhRvnRIu1rbkg6QnZdijciIfY0g3E61+cnO7DD+/UzAuW6JkqL
dchIQuKvcWAtDV9HTakVb/iUQcRSMu11ZZImR/VJqr9zAlV3LsEZ7kKVeL0rqNan
otnDgKb5aNGYkQvX+4gtdzVDxHMlqS2U4s6a58HADO7MFmoa/dBFyg5BEXSSMH9E
V2fwydk3N4sAu79o6osdfIe3Uz6lLk1G0kAJjAoDldu2HGKg1hbNmoMSErLWorL/
B8bWe+gzKIZ9zxAGiU7AuMNdmtnTZcA+kLRoCfmQBAACIqil7SXxHh+LhvfP86V/
h53VHbUBkJv+JoyhiUaMjhJYIT1/BVKOIbWL/HeGpfnY1txmB4+TfF0PsKBro1qv
xrBhUSHynPoiXeJBxVpXZUIrP2q3PSRpVcD7j4k/f5J9ZylMzK1wuaWU96Tu8ve8
5JzHwOzUnHMcucL9q1qGm4Qaq9N9yQTQ3XytEjbAKGY21XtU8vyAEklNxGvP27wm
Kww7c69VBA5m94GbY4dCFdkPWG03rf8ExCFblfXotZm1QNVLfD5IZo2cfmANWqt6
5CMUlhSXF10XljqaWcu8ZEFdzwsj+nO2cyPH+vwCzFPwZznzdynkO1vyMV8P2Wex
Cj53JjQNr/bm7gdSdrZQi+O0Y8clhpgcAc0NH+il0T4OIJ5Tn832OUvOwIiJxRS3
7inmMkC0LY7O56iL05VHmf2i2/JxqjWgH2GonB1QW6OF7dNZvdRN3ZyYQd9hP8Iu
gHuAA7/GewjBTFwCqW+wsHDbsxg26l8KX3WT7NfdlXoNZLxSOThMC0WPTnbrQBKl
FnZ4ttfzTnteSMNRtmnqgcRjRMOOHf6wWYq91AaZfOB9N6ZWexDtOI0Y3Vu2IhZR
uI5QGDwHGNzECSTDxFcMqZNKMazMdSfssH6ANZ/5tzcp6hBgLurhdGEBYaDVpGHg
F3XH/VxjVQro5bfP0F0ANWebojSuO818KKHPGSXma6rLLQ1Nkb2gKH87SRp/H6Ee
KwRosTvx1BKbM3gEZTkP0xmfLA5weAV+GGGxM4YC3LONT7oXmQLtcTODeQ5nY/DS
eaulCK9D8183expDwqPSDxCcJcD6tvpuT0FK6LVuqRo5hXSq7y2fK7Qt2jxNze8W
Rzq8oUoGT46nhFN+a1b2kjg8+zusAdBVt81PFDtnBmpAixekp8vvf3moVlqMmlKo
aCULwE71SKjpGP6Dk3KdZKkIVibOiXJvetOjSRU3KC9L9bDbeJ0lV2Zze7FNM34t
HofJWi1ALlQ0Bm4+xwqm0ut5QkMY8OJZgb70qM0/oBvkOzrJOF+iZuPonp9hErfq
clEvpwisLvjc88qY8E1+n7p7q+UtAq7YZZ700sXLJ94NeKk/nrpxQuhOIUB75k/0
Jh0xVxE6wtZjrSybxJfqHDZzASGwownvTzwjWBJElDghUxOtC3AONy41MoKbTluS
JmN97COMt6EmCbFadg6dUKhQyS8Bm7RboaF9Xhp5ROi4twMyus1l1i973h8aq7VH
KB3ujW7oTuAH4b/q8iwqOxZiK5XspGgNCbXozfS2rnHd99rdCG6lMq+DXWXEhtLA
ly6ckrxVWon8vXM1sYDXZYwrpIOh+hIrIoiN7VrQp3pEepnlUYHtdgMkWVeqeBFW
7NnlSFvTGCvQIl4I0X71EVHaagBOe0yb1NdoJASdofs9xj7A/vq2U0MEersmwJAW
otMltYvJ7fkYJNwFB8qMOenMXEGxYVDDKGC76GZOC54CCv3diDvwzDKJRYoE8zb5
gUwlHLemPLt5mJrgT4jL+7RzE9/f+LwD1HcTrA4YzRv08oJQDY3MZ8sha2aSVKlU
wc19kSPvguqeynnat7r9Wm8NfT5apDVQ7MgyDL3ra8AI7MwheMpf0LhVQJJr4nQX
uccKZ9DepnzcZWfL9FhfLvM/k0ony6a6hSAJRBpKhUsPOOZceiTLdftZekZ5Nu9O
CHTH55GMU9138mhUebcPeejAsNOo9XBWxijm9tO427pjeirU9sO/bhq7wgG81dOC
aTH4ftjZSjyLtSNGz0NXFK4HB9EZ10Il1qZeGmr1U3BYaXHWK404oTxVQ/OCspXf
YLSxg1v/8HHpUaN1/HmICHbri2TJkjn4e50ROhXQ/d+79xycS4gFnh/tzJUMOcs7
j8qsUXJI4qrBdWhkgBoufqH8rvqA+aUnQZKtKYvx5E8riD13K2rtdE5GpoVt8iAd
MfYXgWgZGbJ7BNydEBMNCiRCAPKutcly6TXdbur6LQJOjrpsmzo+cVBFT9+HC81d
hIrQUqRYwGmWJnyLGKhe8rgrYcGVWRArQwJ2V173skxTeLs81YqefcC2xdvoxHjt
GGCJj21C5ixKcpZsUoLKXkoBuTU3urOXEDw5B6QOyWkssGDpgMRH1euLQPbHuOqx
ObFVF6iGlKF77KhunRaMWGpKlbcbXMhqSDmWJFHLNyDTqx0obJG9TIzYk7AqEMEV
VcddF2BYBTY04cIGcHTFE0SAKFBMdQSr0sWLMRGz4TD1xjAVLjZdOEBdwn51jwZz
kIP4GHszoOHbSWZY5UUK5jlNSpBkFDurRjgwrZP8v5wgsAiXdwiqOrg7Ez7dLFFt
3UfZdegjtFdJCczpCU4eVIBCqbUqonznXtQYm8jqb+flr4+KJsWSv0ezJwqIGTQM
z63z8GuIcX+OWvmRb8D4V78HYLyAJQGvHX1IWem4m4UMH0XbIoGv0Zv81s0qLJRm
QOVXhvzvU3HT3KevkysACkdJFBrze4m7/NfYTTABCQoq8EnOgQeKMtcaLgZfZ8LL
Cks7w/M8L9XHvQYoAMPhaojksQvIQoxW8omaTreYYRBYOHnC3FrshWosSy0NGMtz
s5nZGKJxklRofdoNldAYb2kni0jd1HXvJfo2GeQSQwFdqTOD7VDxxZzSUKfHNht+
MPrai7n5hoMZ9lBe+KaobcGVBv7iMFuQh8GjBXCfJDPVsvlj/Fhh7fvKQu0Uh1aL
6/1ICJSt2QN4L0sZ/ETbloopuRdiOm+YcGUS1GCoOdeKFa7G1qDdQq+wzbvYB1qS
YM45Y1J30t1s18wIG0KvariutO8X+zDNtSw80CoHfwEs3EMaqZxsmiCCcJaylN1p
GNMHpbMFDx2v3jt1XHYLUnuWitBeGKlFkTFeDlef6QkhRDvFuBRPeo6i7ajVTinu
9Tr4mdkedR6EfAIacfl1xzTP8fx8joWSzb2b90glS4Bum4vXVxXG1jOVsvcCDt/E
E7oe1GItKVTX/MP40U09Mt97gUM07BqTPoVbHZaZQ5CWLX74uyZggs7aY0tPw0AB
Ot3PIkmU5bq3S/qfyem8Tp3/H7NNpnurrHnGjDKSKELnOIoHt4N+duz8zQHmisBH
cCheRMl+LGmUqqSsonxuGyaFS31wFtrpiPvf5Zg0D6tl71kMiePF1Nh1wB/owR70
s2tycgAfQVP0xcLI5bgBLiOkbdS5tNzdP76ptfhDCHGlCXxxshtEpCa/ycj4r7Pb
Sq1azKDcZbtVCvnqxgX8EMHSf1MczHVOgROoVDbaYUQx+iIjgjdSzmns0mAdDlxf
bgwqu1c/emc+Q2m+ebgItY4wt7zGUYE0MFVX2MP4NSF1SvgfIfE7xLL58GQQnB5p
k4vCLLuFTK/m08VjuKStYGOL8vLzaG7TyELChmIgPiiIRV/o6Bse8pPFfrsOHxs1
IbnK2QRDp91Iz/YYMfRkhmNH+ArN8DN5mx4nuUpNuItVEVsCspdShFWFUZUqeQf9
p2XSKCN2GijZ/8rD9jxkg99AIRE8PJwnaiTr2MdmPL4RSVKomBIhlQNqY3eUtqRK
w04B1s/mi3Udy0pbwTIH8MhCIrAga7Im3qx8zm0q/3A/T/AtZR0HbbFWWdi1jz98
z/bE1qD6WV2jwhZyj7fnljCgAA5oujz1BHADe2pID2z+ksfwtNt+MMlhMgKuRfAB
art4q5D80n5IrA1wrgQFdibQPta2xYlNQPJfEDoeD5OJZ+6cVdwiTwCNuratm4K3
fHNpswjUirvBHya139zjqI3faCGCmGsP8woTyF/asQDIBH/6aNA/cusf34jhH2DX
C9NzeLRfXgkMfEzz2NRCxgmIvw36uoaNVc9KBkm5RdjHGpC9V9QOtqY5hBiVg1i/
OkSk7r2/lnwtAfUfV6i8MvmdoTzl4mFlxrihSD7oVDHwF/+h2cozDSvJ3XGS9z1Z
RAKbxxJ4VX4V8G2Ckz6Aa2N98WEc2gBaY+m+QM0OceexmwXXsun8HhWMaDSTPkjf
tUY9xnBQY413e1LM5PCO6SXrjBPb4YIPEH0GlyQbmQCk8IB0NFC9aiuIK4s2W/sS
k52i0FP6/LhToD9N6kDQWb9qepTn4m6xPAxw7Qz0YmmckNjIujKcHOA1CoD5JWll
o2hoABN0rIfRzdbceUDqgBotDDHzzA+V9IoU50/ueBIqc0omxqGJAg2fInuUSfsG
wKfVqn6NFpYqdhMc+Z+SQkyA6hyG5xnbcdENVNnNMI05gzFjRP40riKhmu8z0GlF
S5/uR9L1awtU1vZSCs4IODBySePLfE1WWNPzup+5E8//N6bAfeObujN8wY4ZW1If
FlB0GB7uJ5YHJi3iRdNimjO6qiYIfQpFO0l65LbO+HL8q2fTM0a0ZGhgc0rCOA8F
KXf/OoLCfwBZysxOUznLSawza67qdqOq1SFpb+GJ4PcIncf7rT7RDGgPkOm1wVXF
WmRhYRX6Qa68KjavsZusG7zDsBvVQ1Jijr1M3cMGvfS+feb4kWyYCFnwmy1Dh1Vw
ksJLDzyzDAkgW4/ayQPZGj7EsW5AIVRXPtRLyhIaYxVnRF69K8A0zZgLRk2gYNV3
Xl8Nx3ew3naLfWOoc9CZzZaiAbM2Z76u7GWTxBrBjuEBgXs4i0qgOMTUC1owP9kq
HJAbhkVTLzPCxfV7b7Do4lqTfyFaCCctvUbfAfLwQXxA9q53FFq97wzcHRsV4ZyK
0VjpprfRLfF54MSYTkYa29mMKsXFrMYOZ+xBuBrO7E7/kmvWnk1iHw9InTD6u81T
NL2KqSWEqjdOlEV8heQId+28bUp/1nGIQa8qAu3zJfC0kZdOKzC20lZNCwqHC++F
/qXJK4oGeLbKbc49AO/N+7QcOb+8lBaNLyBAY5yCv67YGb/Cyg8dWcFwtxTJ5tZf
8vHFCFTzR7wNKjkONZNQTcJpvmvtuwU/MnyYp4pgh03Qak5rkeijotOSH24GnG5F
8fHxc7o9tmk2NmDAdmht2aJmM0aXCdhIENu1wAUxTTuY765RY6Y3ySQOuV07efu6
4TziZ4BFcJZCUwrzoFSAnVoEHPdtAoBMdBuIfXUvzqoijv8E/XKajkfEV02YcXmO
vXUQsEjNakGIY8TLSiPqFBBMgguXI8Xzbv5tRGuDakfdkoTTRxAEU8Psz9C/+4Zh
mo6JuUIvPQjQrGHcS4pDPmMDS5xxKJ4j8thMAvF7ZnqXpDzCix65Q7sACFLJKaEC
OH/3Oub2k9YyO7xC1vdjwxvFccuZoVxpa28qK3p4/HykucssEszDzgTOOI+WOiss
w8zDb7DFH6GZvDuiHlfI5eF/15WaK1kZf6Nf2Kec2UymEJyga2/QtthOacLfcU1d
6HNsTK48L4qCuh86NKscYwJdX4F6zHOmJ364BJWFRUrnagX+fFT0ENzp6Vc4d0/c
3Ehp6NYUcp7kfL/FATP/nmaqKWgoMUuuOC7TYBeD/mhx6CpR9npg+fJyeuLPUSs9
u3v5aNxzZZVHB8bfSwGKNHuWCzfgTpkSJDC3PDaoIb4jYkdvGU9JPzfP5PUI/2PX
f0LeXZQGciY5YNkZFF7MjGtcO8whgzw65phHS2QDe+zcdAn104+2Z5UWT0X7N1ml
ermruvZ7XpMaeLMahdEiVz2/BBCMDSTyAk5kEFcuWl9xx37p+XwxOEvdZah8+4Bo
h9rM/WA3ZB3h54fvYoYOrwtu4nIhbDEISCKCuANzl6xXYs2G0f3vI7Lw+VJIr/Un
IikEa56rxStDKLjLYZIgGQrgCSU+5xU4P6FSM763sXcHQiCpcJ+OGcurgEQRjRRd
w9/hC+KACc+1jKW1ZwKGsY+4pyyWfkeetP72fiGePA0iakO3pIa0KZDVm8AVb12w
4KH/mbSlJ5wbSqDc+sMwno2JwEIwPOEJEujIlz+Op0Fw18J89P41l7SchqGLLlRk
4+cpa4i66YPAB8b8mZhwdEEnlpmRdsLX1u2TnDCW+nHM4EcqC/KiLePo/PHKoZAX
Ld161kMhVNGgOS9ZjfmwkZRTroaekYhAXugWX/H47giaA/OKSWjA6Eap+FoAPBII
kvHN3wfilVhuE3Ls5f4h/7oyQzVWmQMqsD4VCdTSyq1slLfanja7S16gt2DX+Jzo
SKeRootbu4d5/kfaiBCBA0dBOwtR/qstfXvN1ruiNs3OuB7ogfOiBYaC5C8MJAyY
lKhRPCU8bqSFJRcQQ25DjbTVj1wuJKf/6SZeqo0GbFG/ahtVCzzIXH1XiX2J9YvV
GMkW6N/pQ8yflBYrSku9AYov7rPWzU/hltnLvZ3ZDblJ6p8WCohOdFw1zJTbid9c
p6CKa5gmcGY0Pq6j2QPW1NNgulnivD+whSzf+Q7Xk9RffkZdbHjYjo0YF6kXtYM2
lcTj5J11uirlbCQ7XV7/dWRyMZm3dGS1EAuhSBHCIQHPfz1v5L4tMjFVZ9u2t8ax
om09wtNaeucvwfA5VSzLP9WD3Qnt0qNAJ4SBOD5oFXlkuSf7XiZa7Vd5KqNVWFUh
W1tek3amg+C18tfCl85r0GQFVxErw9AU46i67MWiRYOFMmsti5erXTv1eoWd8L+R
p5G0vfyIidUbmu9l53ug564xjSv4E/OymxwqNtBqhgw5b4NkqXojZSiMjX7nZ2al
zFr2au0JX0sAZGPDAFL/4CZuPfWbC6PNBNSsXXoENl721U4VhdN8qkaYkg9lcLoS
yrMa23FwK9QgKl1lpH/WPe+zm4B+TdvKob9xGgrzf8TmEhVuMeBFuOxeXmrOyydY
v06wvAbFQtFE94kr08rKxxczu5NTdj8I/fFGWZPj5VdhfOi+cZ1E1T0UovicVR7K
+NyeRLrUilvnJzead6I/eH/4LQbEdA60w6IYKlJjAG/pK5d0J7tscNpambCqUagA
JfJwCfiRt6yMVd8c7My8faoUCIBf/Fi76gYcjMoq6QUz76QqCNZU5R5EdWaSOT8c
Bn6dBmDy22Dueoi+lpBc9WN3TYJwrdgk1RJK3VtfDTMwbgGHg9DO+lFxgamiGM5X
qGaWcHYORGFKwqWCmFmbO9gO8EbTgFxEkFp0QIDBwrCTXw2jfllcG0ydHM2ktgqJ
Q+oM7bx0EchkuoQFkmGetW/GlwLsNy/QtHojKRFWo/Rwx+RWkDb7017e/oEVAkkV
gFV/CWlFxVketioDjNcWyL6tMWRPjPozpxJ2AmsOArNREfpg60uEYf675AxOSZog
gezeFMMOcHv/jPa4mmqFOdxN0cG0VbW1vLYC4S1Ycc89pzi5YyhcxtYMIbW8Y7o4
G9uXqY487di+yj9kEBDaYzGug/N11AtQQiry85N2pIAbNSsGRcsQIlsZza350YCv
THvIJsZgIPkAwMVOVNQxFI5QxVkkTQNG/bMTKByIptiCiDsVFGVp22qMXp9mt6vX
s25kdlBLcDV6gUePbEQISyWFZJ00EdFOjibkVvLleyflxQFd6fCv4OxIDgXCNhaJ
FvPb7tposvGR8YFjflZ8daqsSsKXG81Bu+0FJ1Ve34akXJTOThfz/Xqro5hX2icD
RSA83Ua36XavrWxUBCfNAjga5WO2K1qM0uMHv7zaz8aZuPrHlYAI7dVKYmMaJQov
wDUGd4CoPjNHvl5y9d/Zeya920Gvd1LSPGOz9bbwpf+bRjX/E4RP2bBmOOKsV8QQ
XRpx6YIjssKMhpsiAB68HrjFYjykCJWJRnxxMmAQg47JN9H5yT05O/kCmTnPhREh
ANKWtDBZGF66MU7dm7pLVHcZ1Cn5CgvwV8wYh9eUwBsKNiBhR6ICCjaTN4Soue/V
uyG0uP//XMwddzn/diWaKUfS+OLCioqJF4DNr/4HgEgvcJcFOpaPngjyWCbixO4T
tXFl3JysL/B+EizVNbzKYe/vItHjHHL1DQ7nIzj3q69ebG6nfEZ3If2X8Hj2kBNw
+fW7hqXY9von78reN9u4ij2liUJvaO4gAU6NVyXOp+binxGB9bQ8x6r4zAGcsv7L
zOonYY13uCRZ6JmyAVgR+SlyAs+MeP6YlpIFtkdOhO/j3mOrpYqF20VhtfYu73qq
EnR6DaKEpxH9Oedqj9vn2OBQ48rBzDwHmBo3H/5pfamPcn84AbYmuSyh6/rK0mXT
pluOtjaJZ7cws+R+9azsctsHBJi/OtxZTdPfxJ6ws1ZJwhts83aOVUhKYTYfSHUz
xLFInuF4/08xw3r9DuJC2dhinhRqlVpOaAb/PI7pMHlpUtA84tpf9F73zNNTUMs2
R+wQ3b0JCjMWfAAKUUKK5zcIjiv7883BV2kFlZuL1XJb0xzPbZtHUuZZPUGarAOM
iU6+ozgHWiBDTyQDUnZHHWOotIeM3PVWA64g3kAPjYupYhBFahC66ZgcGhb/MiZT
nL9DVIGKkBXQQ4jHfD8wUBjpOp2QNwC732kibA3LvROK64imzQcAaXfurNLUIPf2
hQXWCyTbePE7E6frws5JtX8vw1rAM4/tPhx6Kzg7UsiYCsc+ely18Ce9Q5AT1tm1
vCzoEHk27BJ1T7RdMc8P80T+ktp284hI4UgjUByzOXbpNTyBJa5n/mLIHnHtNTV4
ygIrwo72rN/NBBGC9E5mV9Duk+t+osXgLRNBh7g/gy36Xhqx3GWLZ2dU2eteBQbt
JiB6DYeBDXFMLxnWg2QvEYnwrsOfBtGz9SeXx7giPPEiFhPFGO3MRgUZzG4aaCYs
ufUeCdXr+eo7DI16XDeXQRFetV0cSDacMdB3s25rQ///3GmGSNX8XDaOKmAVpH+i
8PKmXiFjgqyG1rmI/OH59I8yjkfoU0fDhQyIJZ5+8x+i4I0pB2ud7Bk6cHAwUohN
3mTOzmp4qc/iDygdbZygfiJwyYpxznoEQ7QaYFpwa4sOlV8YCb1wIWCxFCqA20De
9PJqIcaaXlkKvpT60c0Wf05wphp3iVw3O4MqoMwso88K5MOZUCeNLLu8CgnqT3dY
hLJA4f1IJJGrTXeKqJZgK6/iqDBdgWe8xP1HQrNUzFCTVeQqg6bhUxbcULd5vlN+
MmRpuvSWlUm11ecasXIl40G65fzJBtUvnzQUgXLcaKEedP4yyY31t79io8hrVZd5
HjCRK9NEVJg1av0hEe3HJTVIH5/dv+b6cd9JxZQdtkH/ds6dXNQl126z/YYqP2YV
BIbNgRo9f05Hz0HZ3XbCJO4e82nRuBEcXw2H/8LFNmoMtP3Wf1Q1MJzgKnIAloYZ
CUtSlfCqVH3TEpWRzUuJJDZV6t8kOzVaHKMVsTYIGWaZjpwgsmnTN1WZQYtQjXin
3WppXE1u3qwJ94pP7mpow4fAjokVi8pRYycsgTmW94xVB3d4VIrQzj2gIsjTg7cs
Mt0nBCFhS5kJsPgZD9MuEOx5fXTRaBxlseE7sT0P3deOAmaXkqzcTI1JA3rarKjd
5nFJ7op0l7Ic/kHSUOiLrxsGSsgSnuOAxerQNO0hjHFiSRu48CSdEP8EBf7l8yI4
g+uyC+6QBWXxwRIbqsVtvN15/G/we4GMbOgWoGPibRr9OkPu9f2sQ65ZfhDySptq
Ny/tt0n0hAP5DutbCakc/OVm23rydQ9KSmHZGNPFSPawX8PyRGF8LDoD9lybwHjL
tCEUBb4Fx84wx4HI70MfsLg5lR1uME8FQypFrd9xfofVWA9LhnX0ZFucTQIA3vBB
MKd1gvuX0wVkfIkyba/iQyBXmZcdzyoOYbX2P4GiC9LMD/455z0mIgqwI3vnXi00
zi76/pybeu5pJtaxmTnUR6mzcuoS6K/wv+1cS+2kJw+J/G+5ixGdh3RFn1g5ZODL
KlmkHsGY/0Ppiek4nW0yZl/FNlIOG/EVTyuA7G0dSwyhyPHsDTbHOBzpei02NCFy
FC5d/AoVotustr8dGvcc2TxJ45sgYH9ZNvs213rVrmNikmHKg+ugbh+cot0wG4qW
hPEe6kFSQ71O+fMKaI/kECh233U36E3djNyHnswE28Ni0qDSdDALdc7M6yMv6gTf
GzcH7RSHvyDrJYnOwcSF76/vcO4eFsXEj4TYfWsw3/F1HZkPJnpvoj60Gypl3O/M
wdmqdpyDyZQM5XDnSczFTm6UIbZUFdwq2fRQql6ed4xUuz2JiSoCPGJ1icKVdasW
9B38HeGlSvw6MmeWIFQmGWglNCAx2XWojCRlwHhX3ChapxV6MWqSjSSHxUFLbM0r
NXG6jMfNDLlI+vxfKEyMwZnucNWOmUM+ynxPcMhGCgngAIJBueWM3e6MeuCoyCpb
Dh7ZCjKozuVuur1jRKrtMHsDxp1UMEbYc5gB2jYe50BW5z5N5uneRzxKeUk/U4uy
WxWkCPQmD/3GDh2KLK3rHuH8QgqKIzlxPWBXysBBYGKJs0AnvbKL/k0V8iHFjgU3
d2yMYhGaqDcVzX8HUjAUuX7vIGYNy/W3Xaf59MWXrDdcyPNpv+VVAAonwrXQyR57
xeEDQo768eNc6fyTqE29IQwxtA7wGj8BWCVmpOp33tt65ZrmMuXVIswMwFQZEY66
TH/+ptZGObbctG8vLf/djK6P/7hIh4c5250CWiWAQtu1covHAc8C7J9GD+pbi1QS
H+rFt4VUTyl4eq6maQmFy/Dk3O4c0bfVVicfob7CkCalgyGTHo1E7qWwifgYGrbq
5gWoCGNLCUj891LW2+3O1kyjEPcZBjJvr0X6JrU0NSknPI/xGmGrYywkv1umboyO
4A3cNvsBg2v4gJ0TPOBIaUpJgoD+vRmzTmRhrHmfv4v582uNmymEpha1Y9GEyb6d
XAwy5fSk5qTMbD9RjZmfPL9jR7xg0OyDqBHtWGT4N16+FEu54bmakmrmhnOLu4uB
ufPiSm01x7gVHxqNPgSUtfm0LDgGHR55ZAWBP+4c1Tuw5blj3LUo3EQozY6Pcbds
0nhBtTIVONo7XFoOsaPfcTgJRkQg4hH5NGV0LZE8AlqnLEks4wC9m7lFeGgoxfUp
c+8talmva8e2v3XHCNagleXsMalm9fxkv7WHjK3Uvjh+WTCGxNKrJvYyNeS8SfDo
VNk2sSPZnlJS7FO9v4X8FTSUfYzPibf1d7QCWdk3QNm5feHZgaIJT/HkNhblY4v8
jSVVVR8WfExuBw9M9bt28RnOebqEea/iOjbz0IO0hiwmbFWTrPPun0zRhT5YSp/4
g7p7fhiu4+YTf+KhnnivzgUdRPEH4hsNWwT4roAeMWkKCg0Dxk+NnTwLpyYeZRt1
+n+72McvN+aoimOktZoGw1rMNUSgUSPdZBtR8lzcehJjV11Bcw682VXwZN1A98sV
IHeYo6rzfXqBesVgwMxxuIOp9vofoaNzSAdtt84hBajiBkTWdT9+JpvxY5TlpXoY
S1Dk2sLdqRhkOhOASfOwjOWvYZtVZju4iGr0eOaWU7NhvXzqVHGgOxZRssDqnXot
BIWsU9/FEhjdIhCkdi0Xcq15GV3SIdoZ/Ek3hQdv/g/jmsoe7trFCx0CsKVsd70x
6TmiQkoKxkmT+GVws9s/G/qjnqNasSXtmZdY6sk+Qs6X0Wi4xhKLSJVuYzAqB2YR
kjvdChJ+loeizONEb3t4eLHpT1qYjd9fAQrEELYrGAvnAxjtj2GMPOW2BLHVYsWG
0LkmTZdMenyFYex6mMdeCOtdTE/H2HxAxyLnCLfFCbCBXGQbUNaPknDx2lJnznZD
rlxF0iJv9dYXYriRAU9INybkTJoGMjHu/tenB6LJp0sYhc5UQDX/kWN2s9D5cQDf
0AS0nKa+sVypmsV1eZ/2anJOxAZBbWYChBSNq6Mg6zYuaIuxisWEnp0tHhFLD32S
IjjJR8J6fTRJ7Di4KNQgtbPA50erLse3FPjcBvOjSEtt92QTE1hukBjhttDWMTud
1M1L3I8hMbwuijWJZuGXCnmMskflhM68g4x5Yh0JcoT7Glm0XYMxIbWBCcXdbl0a
L/q03RunxCbBoxhvUX7tzrJN8U2sF0XTckW+IQHooFe6RADbz5PqIRRoaIz7cB1c
nqipne1RFLf6CrptoP0su5CUEjy2sxjyIL+F/AEYAQxd+hByYs0K9xvejIHY8mWD
JU2kVP2KuAf9PJpaRJS2EB2dzTIttnlF3dZ+xA6uVkrcyPO4hLc0HPHlrKTrTUK0
DhAOi5I2LjTl4EONG/CKKbBj5gYzidTXlUtFYUanAsjLQD8nuGZnO1xX/ryovAjJ
Lth6+keIk8wxZ67u/y/MepgTlTGHT06snDob7xqscCTu6ypDyyhEz0NA01MsDjl5
um7sxbTyYz4Pd6iBUI5iDOia8449VIR7Z8/q1xppjwtjrQZQHbm3Y+BzwDg/4VCw
CaBeyqASBJb5T5jkURhZjZEjnTwSmY2fsU/sAbUvH8HqzVraopib/tXYcGww+bYT
j9dWGiOvyZ6ciCbizC3gQD4VjWl2xC2+DCVloP1QYNcbaPDO491ycxHJpSxpm244
HTWYMozuhrIeBioD4suLQ0DOX0ndr4+SrngDBHJtPtHRcYEO5kuk4JprFyt8zZRK
8pStncDjaWMLn1aIb2w/Upw8lgns0kOENzVEavbNCA7Au352JT8isHQ9rrk903lX
RC7baKOEmSlEHGa/KPtkU+G5hv3GN+PaDJCzdijymc/RSpAEkGyzG76zl0hHgfHg
8f4gTTlu8kgT9KrgapbSUgHI+RXrTARdghR2h85feJh76q6fCbfejhzICLyvc92J
9VZn5vdRiL03JjuSGaA8xTliljf6NjIIUB7bsM/P3sdLKuvB87AcFwAshFzoFKf5
M9rw8rsjorwws43sXqBjjgE5nTHXD7wzgLYpUn8Qde8F1XZYyI1Bm7G7/E9CInpz
imNriqmzpfHpNE7BWCxjIE4KzScH8VbEhvr3q723EasucbtYkdxgQwEHM/tkAPEI
/lIUTv/qhtcbCw0Vi9oyF15Ib8vn/wctG+DNJ2bo/KU0ONpzPauOT7i26m4AKPjO
mn18DISCqtJHqY7EmI2J3GFrj7e6yzILoY4H+IQoC/W9WIfW32tcfROmJ+0uGnyL
Iil8GP0YTVQfqj18Y9vb8Glmph0XzGR69p9LESKwJkifgC7HbvQu3aaltOq38+A3
ewgunP7NjrjDyAWZ3C1BdeaSDKLMR7chYBAGwiwHny5Az1QxUGlExE68WDkQFm41
vDs7UR2nNdx5UCL/X5SIf9GX9WaNb4fiuvGNdEvsd9DMKu+5VEoMZT5f5cXz6Ot/
fJw/5GH6g/bb2NZje2U/hyrEna42yAmNTbTyLc7SQ/7fTcTIhGb4wF0+SbfAgHJD
DLDoKZG9AOD9HsMGSGP4QfUk0lqXVnuBU2EU0+bg41L5S6XTeVQy73xVEHOF0epz
BGk2UklzuGpHEHKPjSkvnY/D99g0d1Mgq8nh7NkNrRWQz7Y4q+h9lqErp+1dYyWy
Ae3hm7+gdFtsxkRDPsxCwlZZyua9ImdzJzNn3yEs1lWT8Nhu4ib+2zvozh7VjfqK
CpjegsqXQx5bGZWyueDzaW3INtm7lbNVDKHPRCdJsh39X7VuOPvKVdYDzc8nbkTz
bs/KF9VhFWTLcBrWwyRATEW5jABcr2KXRGp0xf9IxrW9+LPMsg+snJfVTCOgHaKz
P1UqO9UVQQKoDRAbJ0Hi10pzIOYeXCWYSQyPJcb0uZ5DrjcXG0tIhXNIp6A9FouW
sYxb4wxj4G3hAd+LQMcT3VMf8iQEDlGDGqoQjv2w0vk9Q35rUWpbQXlCD2i9jgGu
G4R1EPwCz+TjN0txMHgRy89WHPJKLyEe4+/oOduXmwhcdSyW/4JvuyUzpowZY7Xi
Nvg+isltUwDL1IkhVkeFGkLlNyigNgkH32q+PG2SykjC2bmwTBN+s8gvwN3iqVAX
lY8W/uSMhZ6lnG8P52HFZFoxhdHSe5Q8DmfKwy4JOe/WVay/J3jeB2qRB3FCjjle
Rjp/bTd7gaQYtuvFINv+OsaF1irnIQyF7XWnT0B/aswpk6+2W9RsGr6B1PbjxjIA
/lzhmcoX1yE3ijKDKjqcnKv/8Dzihw4MS09VEXqFxsshR8MN6I21ZGiTGAn7nBEK
jvdPLo62criFH6WKJvOpILWWW0LfKKJOs4rgplgOnrc6Hp3HkN/ekrei6XXxU4Fn
cyOkFo4h/HlrHjGJAQMvtw5CC4VkamInuICdURn1AW9cWAFdPdm1alOh+Nu05PY9
ajdAu4oZ++pfrpoZVw/wJKLqa8mMJfTf15rbH9jpISxVxarAkGhLT143NrCtYhP1
mcqfB+JCcQzGXk7/lsIDuvdYuVoobcm515o6eAUTNJfHHXeahqzIuEgQHQEOKlsc
AK9dLVVDh4GK7heZ1mBlvGeVplVkLXZXSIQ+gXtH9XaNHr8Us0T7DRtTDtymYZ+x
vzuA1O28kOPGMX2PuMcjeMeSNS4r1s7fJz8gX5aCzGOWnHSig/XjARHJJc+8bw/v
isoyYcU0m0sfc6C8TtK+LmkCwNECGPVajhqXdWMnI93CLmX9IN3SqwOOSgz2atW1
Ju67oC8CqsofvuN517UvzihEQ+xEmZmZj8/SWgnx28xk8QlssVeMFf/NtzE8cjGN
1WcTTaZxwNHaWI10UtFq6gVnlG3VJoXelHee6E8Hg09E47M/VPASOfjLCMc3SzuD
B4MkNhmaQh9BfLkk6oV7AUsFo37jbIoFIFbF13butFdL3HhR23jlgHjsftogz0Eh
PAk5PzxAzFXt/2BcJIi+ufvTJNt67lFljGWObW9Ek3UP+QY4ExdsE/1egzRWbRaG
nEKa9NcK1tvPSyGHaRCezPIJTVUhJZOIe1+4TxcbFe6Y1btQllU4Z7pPCrfOOdPK
VvwnZyHhk0snz1KyptntQJRAKC7oSZLmFnGytdJk8BD7jZjDaU8fIsRanP/X50BH
QHrtZLctsUBX44Tgi+2k1sHBe2J4MML7nXGMxX2f6nFD56wj4Xot8O+wFEqaoFy3
nzYd4+53XaHvSVXSXi02YOtsQKzWMfaqSavVTIdJKirJJM6w9Mu89SBD1Uvjf9p9
CSmKmB4yNAsA0ZqnZHcr4u5LFR8XScFJL2F05XjQ0k44J6MuLJ5VhYhm8+9220kY
vNBfqxlXdL3shozrEUKj0grZJWVbm7AImD8daMA8ABSXFOorTo4DRiMJoR1Xfj4N
bnhLNyNgce2c9GA0ilh7O9qMqamNYBx84NLFSqDJSeCpKBlAkooP4qdTL9BfBySr
Gfg8I7qN9yS9freyYKCE8z00nRbeuPdvjoRQc9hnXhGkgm9Pj1GIlomu1k4hh3Rc
JCy0Mk/CgOkdl6lXlGOovCnf0p3pZjBkb0UYpUBfSDjv+3vpOszE2WBlW0hytg9E
FBO1XDizDZMblB5LpCf4pPMBjIWaigqdp/FvjAQaZFQNxmuQkaUFmnZD1wzlyLhM
HVSR3b6uKl8x+MgDyLIM9eVOGoRxa2YoFjL1D2C5KW1Vva43Ik7QCCvu4AWeQiSb
9IQSkpyfSGBigXyxol55tdy+NP+AF+PLSRuItwsntYmlmt5ek+h0hJKzcwnh6Nl7
Y1FQzF+xKUUYq8C9C1hQ/OLC0NlrUV7JGB/yzfMdh087gMsXHyryphI6dGsYviWx
efuwnwpBuzhz8ytnZMCj67O8cCoYtShjHgu5Kq9RVQ7U19k6+JyIBNYTo6c/HDXP
bDq+62n1qjAoCCYyhmWNUxtFbf1oI8YVbPP3eRwEu2gk6B2TWmqvoqPNXXqaKiNQ
pP3k6iZbjQVJOeByTDqhQs29+ju0ljrFCL4MySn7sWZ0K02Z3vxLHDdHCXnTERLA
pJvD8HJQA39QzCsWi3Sdtgj1q8d2NKfGxpY/IGcGzCa9URovCj8rWUAxFFRLGWZp
iOOHai5adeG8yvIXi0m3BI8/JOp0HeOD3YHE6HFL76g+yl6B5eW6PmVyfrgX/3uw
6l7cL+NiqDJ5fQV4TOrK6t0djVTjr0fCA+D9wae9wZsMJ8XQdGl2+0V7TsLc77bw
sCs18S5Ad+epH+RGtHVtPCiw/098QeO1V9cI8hdAvUaqiBxtT4p1mhbO9U6wxNvB
5FIp4QPIHeQSYIOhHZNJtheU7OpdQnnFHIBtqXUg6rc93Dz1fPNAmt64t+HL/F0U
yeNghhzGSmuRY/ib3U2+74UuhI8EFzXCKX3A+rePjStDTyzX0O9R1bXwbuGUqO9q
aKtXy/wCNHkO5l+uAk5JINEAiS3UWERM6m/Z5IyOcu5Ser2oKiInKyCaS9xGff78
+YL6NyfNWwOmB+p5nlexCw6t1z8+DJ3eFdhexdixy+StBC4govYZEYGQNPDfkD9H
Ai/G5i6yy+JbuoWDnryQ5VQe+u04RJc92EwNRJXpKoMvRyg8cZczKA4Yf7uauY/i
cUvau1kRbwA8vXid2ys7gp2j7w+YjdLkEsnfN6eGb5l/V0DxHFMSU9RNkUS3xpr/
WAfRtd47ubkWQljYUQ0or+oxALB3BptJXRUu0kZSe19EBSHeVOVGO6TbEOw152+o
JDsHmUnsPmnqyho/VLMLjxgUVJtCfLAtZ+8cfomwvaxMLQ3x4Y7t5O7J8l9TIW6N
Ymrk2577rUbcKEZUqkLlBwzm7PNQEGHNZovDTGpE/x74EAMxMpxeowITWZDwxwWD
6AVc6q2ARXlhcyif5IFfuJbsSPZtAgnU+bM2001xA3BCaf3vIBtmo1uiRSS5hlPU
t6K2acn1e9QZ9vmg3ZgVL8+7Uk3A55W6zoBsCfbKNXUh0fH1p9bSc7s58vQWr4T5
L48sg6lPu/n3vArwYrO49kunQS0iGSG4P6yI+9KrNZQhhwIV8XBBWosn7PevBi4c
4/WueuXHAL/TF9DoSzHTgQ1sITF/5/1KsJ+u9IGlvGoItpyvr+yWK7jZaWcSoNUI
qnoWpVu+P9+VZQXiViibD6+GxhBgV7CiFN9Kam9s+lLCj8rMXkZCPLJXdBlNndv8
7sQo50hJ0nVI/Z8wTbjF5JenOZ13kbJD5RIovib1nIm4oJEfsTLCh+6yhu+m9hoi
eOw0gYbxUgkYqZO2l1hYZ7rzfS5yLz4Dq+/uvyZrx5lwYHlwEAZWCSj9DbsaQe0I
6xmA0mgqsf6fyln7JtY5VCex2n4QoL4oB0e3Z6qvueMiNrPfZhUgKzeq2/ZA+fTW
Uf7dk7pqXsqQ28eB597+gWUQzraWP5XfD+Mn5G79gye0xdq7OeE0GhRpP536F6CN
qvqrcr3OwLf45UV4S+SSJGXf6YyS0XK2CSptg/+zuSKwJXoiJS9nsNoOzLUjCx2T
yAtYEdBaEOofbfAwvhqOE72ud2a2I8UCBTFl1OgpkVT6c7DROBpgHxzHph+pwLtf
kmUxVXIbU+/MCvC+H1HghQe97aEZFSE8bKjDWoIOJXP3Tt25onQHzrizgMV7wRMW
uB3WiToZkWMnkz7OcjRajsDzT6CuKjNnwTsV7wEoAI45Quv3SW/tgdZPH0KzCyPv
pZHCZ68rNWMCxvDQbKZujKzkUaLyMzPkh7GUL14VQMaWAbQovC3BDY/kGBsBy53F
P9BGQ10Wev1ti7GokpDtHKvfDtUHN2FOtZgd1GhY2MSRttnWsFkbBvphjYo+LKO0
234BV1enEfPeYl+R37QDwTz3zD64EgJ2QB+sIg17kIYR8saMzSXZ5zl71IOM3Vma
YdtiYYjT/Wav4hUtZIw/W4k2JaRCoq8q4sprxBZ1fAk6xMHCPMOITu/0qVXJllIn
N+8WMhW1G6o4sNlDvwHGgzWuKO+bDmZPyQdOXHQ6RjC5wi9q3sUYzDPxUcdU6JUz
oOvPNnoi0RhcW2uSw5RyBXKWCQAfRoCQZ/Oqx5pBRkysMloIXFBMq7OLzB4r0QQ7
KQnrlmzSMtmpcvW9efmUNVqs8IVJJK3qTxWnrndRsi7RbKVcOGeohsSOcbJmbD9g
3XTIlpZonIVaGRHyynBd6AslXDqLyQljnAVYJJD12Z/KTCnbVyx3zUi+ytOqfbrm
tRUtpuxtt6JiMmcE5R7DZxUbhRWdwTggKBDE5cCK/G3gsSWyWLByawuDq5FNS4wr
FPaN+iH2Z+eqC38ptZkwOZRtlDf+495oE/Cw6s6LpNj/4hru1z+c+teFP7HN+UIh
yklRsSUHErg7YhgZT5roYfOarH04wqqAlebdeEioTUGPJDufsT5HGoW4LMtc8PgE
WtZrW1HpVE3Tnn4jUYShsFtfPEY0N6Lf7iztq5wvXceapTmH0Q7BUKOVfrEPCbxu
jEuSmmIW1z8xT3QfusuJKtu39BpvkxW5IFogDduROTFgTOTnW66LTa9+X5WGDomu
QYDYZMPp8WdU/bA2rWJetDVpKsKhe2Fo/QAgG/XRYZDsprCoebRhjC1sgfiqsCTq
n8qS+kgNk+m1z79cK1WwNuiVgZQMqa1XnMOWGIuB8u/lJrckZnYVg10kmfuisGgg
ZtPtj2NssU+H4Twe4KTXjBcr1hapzfKa6uRpdAqk4FMP1UXwQUoFeHSPXKPH6gtv
/dj1XbGsWxpglu0xZenW/Z3JV+emZSVlVu4bvP4leuKZWRtQIQBuBEbD+f+ZaFj/
HBn3VY8UawJVlVwwZ6LIuoh+zPuvRjVprT+SstSmRY+4zCwKY5vr8CXAcBVFlXtX
X50FXje/Yw5BNzJvgi7ZzZaoc0R+b2bqC5+oJFrbDaKDTLXnCaiDaQJT5+Nkepj/
NnL371roTRo6tGcEDxNo5+fSaprnEMhkwPeyKaTH3TB229pyP1Dy4p1l/lyNzbp0
jx4wGeirprsLAiDBY5TlYy/b+b7IEKccH4bvlGV8dMCQubAL/MxkKbtn5t4of24+
czaEgG6Wn3cH434/j85D2OvXZQM/OtxQxH7x7hl3nCA9wcqaECdc2NLjf7MQtC10
1HLNJMqkG667z4JWmiomKB9C1tzoPjp1/M5ao1fbFAdK+vMQm6SvbB7SzkdkxkA8
ApAdcfSQxrEDvLQT8JpMzfo4dNrlISOT5PBWMqxPcklLvjmOjAU2GuuuE2Ma1ZYQ
/olJpdDUfVOKgOSaiAHixMrTVHCtsfpKuoI/DXF5UKiROSuesV3sM1IoCs8lz2HL
D0p7v+ZxmLV8fbVw22yQlVGNlddDqRsRqfzW2OkQ6NWiQEaTAuBj8gFxmjn1Qjrx
u7ElUfTHLEq/htDiDY234FEGUtSlI02f+sSsuYIJF4aGE6urIHIgSU9lHaH39hX3
CljMMaExKppqO1GL9cYOzyvi/ouxCSX12pbKd5/YgpzVUj3ki/uXnNgnD/YnG6J4
DaYXi9HPTM95K31P0cIPFEKfVdRiPZrbxZxaNLKRy5o2tcZZJDS8dpp1h7ZYkH/4
GQaRRNZ8VN+igaaE/jGJLGNFeAdyGTMy7fTUuYfPlwx3zRSiB5vPVwFyus5yPB8y
2J3od03oJAzcI1I0F5O1nVDThFZz8iHNwcNZ/FWWCScxAAK3HAiczSLIqJ4aFv7o
Xsmnv0bXr9z2hBHiqZdHpWkGTdKLyKX3GOKt2xEn/xR8BoBOG7lFzRpotAqIr6Kn
N7VVlEtY/UugnREXST4z3uNxWQ/iImchKvxwxpuuhIX2paNgmfdQ+c5hhUnAQbYk
V93pzMRg9Uyx3OBS3ZWOij9H9Y4UuWzUGpNrXDpJxPT9XnuRxuOjb5wN9ra4oGdt
S26Ex1c5mkTCpihz/LrCNHm+ca+YBSze45m+CXh5qZqtKy1Cp0iyoMYO4mreNodj
ZdAeWsNRdw0wxXghf+gEi19O0c4iA6ZVdt44qQD0Da824Wegn8T2pERIEHADbmJo
hG2w8HuOFUhtdtUhN+p4XxN6w44xFSS829j+AC/Fe677R8zmA9Cr/53JJWOudJBd
2EarEs+GJUukkcXJTqUGujTI7ymkd3+cWON8PWR+RPHIHpWQnGWIArD3EwEUQ8Zi
Q1RSuhedxkXyEeGVZZimmp+WVtkNowYULJ1xEC+6tfGWBPhMOfgK4e+O3qRwBU8F
Y1nZOgsQLdWXnH5nXNYkDx4a52upccI0KU45k+QCCIY5e19HZxlirG6IAK55w4TC
YlBbYodXzchtPytWpvDRYUFSyPhsboaPrZ7i7h4tOb3UoVZVi9Z6KuYGlvc6ppvi
UisTCrBTYSU/5Kds6h+wfKUgu1shaTlCLsLVtQTZEOtZmNx2qyaogBUfxm9NUsrT
Ya83P/3Xj0n1c7hsgf6FVB8WrgBV7oB5OCi4GxFVJfiRlWaKp4vHi8pzVxq2H6DM
M3rkZCyAnKKfqn6JMEGum8/MdpUGsCadCJUPEdF3PRJ6bSgWuq1UG30KplJL61ua
xx+BqhICV1WS/B0KDQ61116QfPc4bihHxDHbP0KRbRuTXcPLPjw8+87PXFpK2YKp
zkjW0qY5NrRX8gnjhnRIpThf4F6iLQ4A2q36ZQrOipaLfxhEvCVWdFYAUYUPjnUr
v7PtGhANyHc12o+20Cth9gcyVHHqVJxGgUebisGIZY1loTmx71n79uS0IY3C83zI
Sl2t5Doy2y593dgr7B5j8WPNacrnZvlVk2A5SZt238DybhXK2u0tfMhDThz15Irp
hNvkJ6gV045PGs+lj0OZ5el0D6o46/VDMw2CbY5DQhQQTFfYmFh6+ZFRyCj47JOr
RAwrrM5pYWH9DGD0qwQ+nsFXR0w1WbgZWUgZXLq/VF6z5hY5Lw+f28Fm4jq9s8Pr
vKDw2z50npQSrQ3Mff+A3VgZcWacpLo+1ImYMkz07HhSd1nCo3GLWBawiC8/tijX
e4hzwue7pktzSzvGP8DHXL2DMKZEoOgSl20XDaqDHdBDRqD+gueZWbZ4pTPK6cop
XTQPM+N6e4IYI123udFo6faUsRdKoYK7e7KiDgkiuo/HuJcGWUhA85S8FKA4l0FM
vda/DgcO8yEcGS3lcDXww+K6zLyE8+0/AMQ3IjG/jIzBYio84SNwxf+KM1nr3f3m
Ek2ZAu1QJDq5FPSox7rrakesHTIeoxtqGavO2WhLhG2/yi3A+nslMZ6bofJGjwn2
4Pp0n6HK0W7SXWAnBJs3LdANpIaRl79mV4LVo559swApFdazNVRDegwbnDZeBjEy
EA8Mdk1L2nsYrbd5Jmx2tAtEnjsgfxdDURogYg3o7TYkTgTWH76pruQyPDi/83Qe
nmaEMFIK0o3X0AsveW4g6KikZeSSqJcrOxib3YdSsYoifFrttaezzCNhQOHeptQ8
L+3ETtrOimI6wK5asp299T324ergTSZEC6ZipjiZgl/ZOse/XRGuDdCAEIwS3NWF
JS0CqZU8HLmKj2nG8XVm46L02HBk/lt+giOZcqQban6vFjCKyO37vUBkgGVSkQbK
PT4wpVgc4wQTry8ah9A09mwZt8EUIpuy6MmSy/TDT7WmiEOH4heMFbuV7HO2jii/
GPNxvBhgfxPFYr4wN0z07oAgXf9cET4/rfmp1YpQljLp2WGjKaiOyg1PCAvDNroT
acoBC1OFU5yqopBjMVH5msssiQZuJbarr5Rl4jk44WYqZt5uHFjZq1AS1dyBWcT6
GIOKhEeIq4ECl94jXZPzoszle0/X9vu/vpjOCdPwLCfF/WKMBOJm/ff2ZfrvoVNV
192wfVW/GI8Xq5g0CkUHBJhE1HmqlQFUEgnN6KCbX+fVhVA98r27GtUUmIMunEDz
jJpBH4gRbygKTeny/a9/RZQ+t4jHfUnYV6TezqbJ5jgX59fk5dQ0G/qh4F6/V1rf
txYyiHMnnVnsy0niN+LoNtBzUFx92js+Ck5LyIyWfDglOlfULB67bUTou59a7n2/
mhSxu0txBucCK6znQRDKUBO2fI4LLx4QNNvf60M3U0EegTWdTigE2GiLrIwJqoFQ
SlyslpXsRwvS5BR2j6U3NCu3FOCOssD/y1kZ/IVEZpBXBbYBvqTyxAMdQmHE/mJC
TbYZBVLn2Q7gcmbIKcX9VoKLqCRJ0ljDYVcwJjACGQbFyz3c8/J7Njp9QO57BhUb
Sj/rNFgYIqPXKkHh16ONxkLi5aALEZba8tnMzYMViNm1XiaeysR5aQp7TdjdAKXi
igdNSmWdQImHK2/0nMO8u4UdWhyoUqgMxUsNyr1eGMPo+VoxnWjZnVfpO47VLl8w
6BhfCElgVHVgzilBNhx3Ip5JEE3moGIcRDnJwbbK7eIfUsb7PNCdlhquzHdwQ63S
yEwSKPFSgfCVWZpxIzCeWsJIYFh46Vl10ORqIv+coevxCpIHkK2c8GhowTxZNtXn
h1Py/StFiVZU9JhurcZTwETbpfgjHEyC1c5atGzzQAbLe/Y+3MkpLGMJjLIAV/az
r+bM5Pe+XyJrpfr6rHup3hjI+BnDmphyOwdm4WPicuErQt9YDfeNjib4YB5Bd4pR
wEkO+gR+5fVDIl10SqYZKYLy0XwW7QDq8vhLZ27ehSzKzWeXAHeq1NE2QHoEK21a
D1SPqEZafqG9YcoUy/YiGco7KtpEZ+TfGJw96QlIRgtEWnNSrxcZvzLRKFTfW0IM
ia9TRgVpvhL+h1yIvaiBGodVINc/rxBrjWs70a/dHeFVsLDL5D4PAaUZJivyfMSC
GsWt5B6875BMyaiUjYo+m6IKEgskwFlpWmhLTMzKC5OcpYnosYHqxY+ZwGdhBYET
lKem6coPEugSxNjbVquShL5geU7SlGrPj/33JewT9eEH2Mhb4QwcI4AnN3yS1/mc
+zYb9ilxA/9I2XNLnMgGreZlIk0zrRsqTuINLgqVbdRMrX3kvuHi9NTHZDVbVWFU
NBQj9u6BwTHBSpuFPAc+lzBteRYxcEDM3Kyv4pR2aW1Bl94cdguLJgiOF4fnC2ud
gkb6S+XHPZnnOosv1lWrjTxgPP62osqkruSo9LT4djCp1ddYqf5msCf1YsIAvgQ6
8KQFZjfGDCx7+dyAlDtsaWs9w0EQDubfi54gQjbhsmFo8QVoeRs+VvDc/P91E/ux
G1EJEMlp334nNJLk6p80zVK47te/kSrLZARqzmMEH8SHpBN1MuYqmR5HBneA4lUm
sEThKnn7+lhlOOA8EhZROLV/MtghwaHfUt1FQq9LPzdqR+hLmqTO8czqGgLMa6VE
6TjM2thCWgplrF561jzO3AiVk17C7Uy/f8dkmYGQsCfPfLyDKu8gL02T4y9W4R5g
pjv/3JFU1Fu9roqph/g7YldwF47Kkg3KyIjTtSLZ0c7+1M2dd4yzDhhu4u8zdACd
VEGSHS/EROukZ50cdnx7ArmJETQkmSxGTOP6wPpKXsp8uraEBIQtscuUh6OvOSX1
1d9hgkEwlK9jop7647iu9E8kM5evrqrlFVinH+xRXUS+bHfGcSIUtifV1xl52p/k
0VL9zkJIRdt+gw7gJTBNLUuoqo6uKpaoMAn0QUA7Q1CKevl1QEZ7d3T/I1B9q5cs
ZhLUCZh76057qGLOdoVxt1YDeQcy5EbngPVZJHdMcdeVNm237WKNN8QdzePikrwO
9i98T2H44WGQm5GZs05UDRz7AtwENgiYyJLWiRYZP1mlsNXm0notkpxD0Ky8WGTw
4miu1B7ChLyWLuxok/nHygU9yo656RjMKgtcMSIZVH5+yPxboRmIbwLAJ7XmE27L
UKfNOjKyp5O4GuIC0nQ/p1/MmVQdPoMZbJMEqwEzHyVOONV68boIOP7MTYkQK+jR
v/Rutv+kGTJlJzR1FeRvqMMfM8RqdyNCYrrc47H/TnS3bxnQzE12pl1hAgrKFH9a
8SxvZK72xt/DL/U1ffd0MsqMV21fHiUKVoDJsB9dvAJay+HDTSGgy1QPijIGlVHO
6HtBa3tnQKqggdi8ei2EUh9mbko2swrB/ONDogXjh2kL/mOX/0lQJCt+Un0jQ0iF
oNhbK6nBO3tG+Iv1vst/tdhjY2bSA8BqDt2qTPQrU1MmiMg7bvXUrsHxwsbjAZQr
JzZU3o3VgP7mWlIGwD6BoJvEGHrjn5Id3QemCDE+xbWigC1EOm9A5PAdzOhi+2tt
OtAgvCoGXjDh1jpNXChw2YOjd5XXbFGcm+/NEgtfmFW2alJJ7drpg45POrciVaLD
cheQJKtIkDuZAfGSQca89VVUggf2/X8iiqWFu1jNq1r9eudAb5fk89Sc3u9McOSL
mlvaa2Y8EToNeYTLMW6rjWdehsPEJKt9vefUZ3KwTHjJGFf+4mroOhhEtUloQ0tf
iIIdRWU5IUjNblNsfOMIra0R9kMpnbMNuEwjuG2EyQ9m40OxidIKjWMP5T2z3DWy
Xb/Pv2TP1KclBUFuy7YxZ7IeSV55nhg2DVMFFwwn5PSexOfYssXcOvz7SCzOIJCK
C1KCTctt4hUTU8oG0voYe29DsHbhlB7DNf1asB9IMDt9VccTiSOO1yaPYvzYH8ss
xVPbATe4pX4ha8ea/HaKwRf43suaohaaRJuwM7/7zNuZAOZIvQ18lMEe3n+Mg+HJ
7DXM5dZWn3j8X+r8CKSmSKJZ3qRUUZ1zPrMsK0YbzfYRTdccET0GdyqqSS3swdlL
KGTSfSvUmlKDAtwLPs+kNTleIQ5nQfNP2oX/2NV4TuTKoyK2kj+sIy5TfE7fV9UV
PteIAPJqTT3aMf7EmJB8M8huRQBmAILjfMDRJzGoKbiDq3vNfHV9fSyJ2eK8unxN
3GCvAfRLNaVA+rvLggRlQL302IOjVD6kDE3Pnbyj7vsPHUqNZuFnhYLGdhhCksCW
bQgFfxToRQ3FXyuWQjv+tjza582b1lF9v7CMF38wMVOIMeScyWKGxA5EQaFyD56N
IYk1xMFuWPRHGNzPBiscJH9rkQ8S3XPxNVxr4ZfewrU0pVCvRFhtB2w7Bl+BugSN
vzHpVcm2m4M21XG909nsS6qhGpWQWabiGC8Hf1f9isypqha2w1K7vDwRd7IuVlkk
zh6519g1+/r7lqvAXJUtwy9aTGgWtOqbp5Ywdy27lW7KdgDAFgLnSgOjcaEblXXW
9UERJl0/sawrnctMm2JlXfhQcyvM7RfP0wHqX/fKMeDLYwraAs9g+M5BICFCQGeb
otm5Rxp5AQ35GKXuIK/jlwUjVATsma9sREJcvtjX3f2Yn/C5pjIYKcMlQhYkhCuk
XozZgmwC1rZOSe6YuQrU9l6rCCpryaokSvwKbNGtvc4nwDefTvWd/zUKuPWpUe42
OoRA4CTEybYTLdtqd9agnU77osW5JrE5PD0tMB/LxIjVbfKEzSzp9rlLHFsCpftO
+oqePIo+B6SEV2J6dKdqemUQq0ZzYL6CAeH2ZYvMJsoTgH5PdfyhQbOBZjZi2bOm
k3Vid87SD3e0lddCt4ojojtQdk2RHDxmpLDyUGRi4+XeMhTznb0rE0JBC6DY0Dk8
sdJEC63FdA5nwa1ozpZ8nq4kdzkBhsL68NwnFUij+YvIi7YxFlS6HxDOtqCHWl4v
/Ft/EMot2G7CF7NB1I9T3oP2CinnHnnDgyNuyenDpOdQH+EP/9NOB1gVcISuY+RU
YeZPv74hYF5p/T+NKYH934AIn9665u4esITGZMZ9kunj5fwvYH8rV8mBuJB5ronF
8c8ZmUN2/AasitluEEVdqhZPpCA87MMurNKvo5D6Aa0eRsvg/+pbMJV6CDZQ6P01
FLPs3x0BM/q8myj5Qrg8kFYoyN4ZEoMMVfHdsoW311mhP15kYkA09DfVggW02Bkn
WJasVV9zlZsrdJTgoEUL4Uh39EP3Wi3b7l/D+KGj2OcEsd4QPdRaOEtyWUFuYI8A
sojtLiKqoZVr6UHBsZ/lOva/u1XPiBuU5ZsfWFPinK3YV1++O7N26xTJi44zzWcy
Le0ExeoiqkYvPdMuQRbKukZJSTedt6d7HKwY2h7Qyb30bpPTrGedLAa/GiTqDBve
neKmNNlfMkEnBc7/IQ7X9eVRPlQFMyZQaXCc6qlEyRKX7Z6B3hJhkwe24NZEoVk/
BvooR0jfGta+IaOOm6xxVr/vLBRfxVP3BiKjBm5F/NNtLVW9rjUSBeW4xrzKEcp3
GWeX9ZQTyMZ4TBt6mCxAjNzYCLi2101uJUmbCzpFBEvbWjGGfRT6rbNF+IsUblCJ
Fcdc67KGNvzdclH8CoeqLiEh0EvPOztaf/3mX55QGXoJbzqw/0TWIupGyE40U8zs
NW7WcB0VYTdMI0sxzxa/T3dOR+xYqT/B46CMUvYqClgx70VBYPOwwOs1ccCW2cHf
6O3IUiEgywfDPi9QpmtyAO+oOfiHV3YRFrnPr/aUN9jsqvgOMKwPjjE+nSJxHa9X
VqS9Xvrk3OzYsyLzT6BqqO/VrujF0A+wGxBJI7yBwcYBDBIyw3g24t79YJzfhV7J
3RBtOZIFwGySw3V2Up1gYmd4A2olPleQOPmd+rwNHIBhjCdd2s3zT1PXWwaEiBDS
C0sQxNrw87J8Vled6yt3S6E6xJj8RDbavW8IW5QkpK12v6KZl8+A/5n6LoepchUP
/RihQoAnn/0TynIZ26hBGy01QM0cGNDq/WFRr30XzrfGjCy9JT0m1Pses52kXGNA
8sRBGAxuFHjyq44BjPQGKIG5c1cNG/zyv70+lc9ITgValKJlZI9zNgNfGTBbrpmO
VkgCma1IZkwYk1LI39s/ENmp9Ot+AiULOW/ej5RRJR7lR0yftJSXq1ngqZfSvvjC
Qkuw5NkppAc2eX5jJ95QnUjh/NiA/5s227w8M87VWaW9MWtkpIOCXUeA/NnXca60
LIyryiUhD+KrFUkzW43KhlkNRuHnFJ+RyiPqvaVtYkyZdlQvncXiUfLbjlznFuF+
3MZ1T1orwQ+DmGWoqAloD2JVAJGKbxt6iyotjnGOEr/g2wdv9cEACDrVc9OQNfzq
/QQ3k5modzletjC2vA6S97hB0syFHMqANPYBr3Wpqo3Jx1VX65DM4YTuIpGhxnWz
+f5miAuHsHYLGcXLQYVOBomyt32uEVx40WaiPSdVV4Ybs1tBwixuggbtDNAOw83y
LI1ZM+PWtB+1V5/XnjaQdP44etsoV+Q+W4FoCfCg+FumLVnunVl59oAhNk16nkD4
TYBbkynqcIzuFpvfXg68aQx/2TThbVbKu7UT2Lg4FI9GfsoLL8uhyg5gMBc5W4Ot
oJpAF6PJrytN6yEorR0rBnW7fyRP+QBI1AUgSrsYzTNcdmUd0cs2/u9TcMtECbLj
weORaq69s/qPNK+PiHtuhWYd/Bd23+I4+ikdCkArCR6xA1KHZAptC36vSdSMQ3O0
PUiRZcYxZV+DQ/I7zjKjZ4PI/2zMHW1bfSGNSR77rlmeJEvK7VG8LnuR4LKCC/IM
5rMq3t0xqb7GeZD4XMhN/H3QMocXNfymrRWGsOfvait1LHtc+XG+Kih8jxIb2F78
7tLq09VhneZq5Z6/rqSe7wa4jHI7Iq+j8kquqzwhz3iOM6yPvgTNvsE9LP6WGtJE
WSVwIJ5OUMXkFlUIft9ZzwW6I5yo40CrX0hbygRMDJHBp1YuzeGDBclDfOt59AQ4
yZQYWtOObsz7q+cl7mFUeD5HP/cQxs3Hfcs0yCMDtRor336LzGbSAWCFf/wdgzOS
oxccQ1c7qNhjFy7EvFcig/FxD1c5K+zKuuR9HyQLLZKJ08mp1CI2ojLFvTl1cJ01
Fj1bq96idHaJKcLQeFTycCV1G5wdCmUoEIDnfpM4JWMJa8wry0P5rh9XQxFFmIwj
epYWyAM4bQCQwjeOPrdJoSJvaOdzTIK6PvxUchsazTsIfrKL2X5dZlNGbrbxKpb2
I7s8jDPyvfVA/Q6V5R4A/K4Dgjj3pimtC5+ITLSLOI/vXQPYCF4S2B958J7pQae3
zBOi2PgxGmh63+wTRaq9uEy78UOkYqm9FM3y0UnEUFEFWgJM3wSS5jgTVPStD4OY
cXFPdgsye0qpUvKJYMPJkpPOKVXMeNQrNMLE8A0Jq4e/PFPxCfqB+6llf4gc/OT4
3heeQqPkUapjNlgnQaK0H5Fdr4CmeCrdwkFm5pJBot7Xk+2BIJEJpoV1SyTkayTb
9+oYu2g6eivpZzuGXIKDPtsbsPQlS0/inrgFr9T2yuK17bMUMqBfoibHbzWcjev+
SC7t7EE5zVZUWexCTL2nTlYAZ09iCO0hApi6BfAPh6LxQ/yccj/X5RYHPVo5ta+k
t17uh0Y/BeKsNONlpH1d80pyT1G3JTix3q9KIRYzpbIlaIcXV6Iq7I1I+khAjNuK
wzdxEoijgpkWaXtV074/Lw56/Ree0QgaLhlhBCSwlkHuOY5jzGZZb5T8+i1S6WcR
QZoF6i/wmGDPA3t0nuW5ok2Af6YC30qwX57XjDCf5YDmqjp/YHaRvfXMXGpNKs76
w08ff7vxf6CDG4dBkomNAfqM5NBbOaVnFhwOE5ck3sOjHS1OXs/9AYl3n+/DjdDB
IzORZcSxq8WLDzjqsUw6+oQ4t1sX4HrSklt2eRi95ioSu0nqsMvdmArr5BDqgHML
AB87ik52r7GxkhWvFDAbtOD0kxYg5YIqB5/7RbOsQMat00jXGPmPMy8y8DpeibNc
0dmy1ZAbzKd7yo+wdM0lAfUskeb1X7VB8FtUmq39T8iyo5cdrEljrIuppcqlrxTS
ezCtun9mjKDy9tjYuv0fsTW+CAXaKb41phRDraSj37djqlprsPOvLMRXthmFAE1O
yHwAyItfJrPO/x7JhadDeKLVWHwlbMnWUzYdG/oR7ln7YWNDnwOwISUU9WtlzE7f
koHddD/9GPHDytwMfkXKlpxoG+Na4Id/ECtDVThjRnOXIrIMtrqqBnKFZAiS0ARb
0ng+yEkJEDBP9qG5FM/BBfxrJt7+MxiPjYqhdQmVdV5WRXbL1+2sWLlcYzUNGUIn
ghSD80Xyd1FDRqkYd649plq0Kkfj733xpwXB3FuvZsSY34cbU7iYW1BriAYalOdQ
gNVW3x8rDzVCQ4KIdnqzm8uQYLLAgt9hdK5aDQB3l4EeQ1MRxXZMtJTHoVCB8Pk7
dQOq26x22YZQ3lf4zs0tzL8uwRKkvU6cUwPqzC5Quizk0aQBCfkjtn9t9mB06n0B
KArfy/YNmR6WDrY2SVH0hXf321ZDwKPm7OI5JdoCBHximsvv11XxLuUavJu8fzxE
++kORnis2S6UUCwZEdt1wScW44N1gsuqyl2/fqSU0OnFapiS4AjQaLPadxoPU3ju
kcWhU1v/0GreQp/wUK46AOg9O+E165JQwOa9lKaufaLECf7+Gc/KLqk/yaRmpyOP
9qX6vO1vOITOOM5Ue1Teaul7ZuDd6wfXgH09v5XHetFLKU4Q7st3h87I7SHN/RbJ
WG8oRSFPL5yF1FxJRRmLZ6NkOSZMLqe6nDNPbpw7TrtmM+moQxdjH4+ydMh6dU64
0ZTgkOwCjE5vhtY+xSixY88zq+xY5uIx4g4gu52LlNqZwcl84QcYK7aVQkenVUWB
EErbmLy7fsdB+ByoXv110yyEkn09+uVkOSl8tbnXo7TKTVILKlCz2BU3XPrw93CQ
NsxDAL+hvIXCkt6wy06p5AbKxvF0zUwgwOWklDD9qmf0eNjnVb/1gia/C/EnlkFs
lkBNFvSzFZ+p0I5FWljSKcp4F8iyEILa4PNiI0uvydyefvfxZiSy0J1yHHwHkced
cFzkAYs8MCI4j3QMJ7RpWUXda076IBo2fiBCxFiXJ9nzhUauvX3eHV1PQ8/sZyeb
nfEmm1xdiqNGU7qlZ/Rv4GVDYSMki8tE/fij+a2Jo+l+Mf903gs1ldyVZ0VhPVIy
/FjLQGWAhQaDnJM0DZvsgYqBn+KVYfR09jUK7eHR6YUZTBRf6KQAPVR+nrh9QIjL
JTyu4Gwzt2vs0U5c2DjLSMnf0U5RLnEPtKn1w8sHqXi0SMFIfQc6UnJHaj9HXgpe
wT8KJghcUNPI8laqIGv38PPWqiQNwGOvwTPdoPKoBZn6yoMyIap1aD0QNADZOEXw
C67pJ4FCFQh4yiX4EdmmgmR9I+Vi0niGosYpWgYqJqXlwIz9o4Wsw0r9aGslIabl
X9tJtlzZe+J1BJajUGBY+bR6KE979HZ639+oG4RKcJhZAz9LdXhMF5SOo9Z/sKtj
pq0+qHTqQhM2ZpetiThsMR2v/ABNJQwqa0N9ygFAvj6LMUwU3yKm3WoILFlaJvJl
LgZ5ofdTUpYZSgtFuaf2Q91gJPl+NcWwdgksQ3r+Is4EMvMqmp94gvrvjvGrtWJY
jV1Aj7ePOL7jn5St5GCCgyhVnJDit8UW2ZQw7+pwSHyO74X1E7cRr902D1zofjji
d24Vxe0d1dW1hsagpwlO7N9FpZLt5+xbi3l+pZ85xPPC7YavTMVlPQgwmxEz7dPl
gFE41ewEgQNTvPEV3saC6PJ8yrxsmbPodI8FxECA8tOyHJH2EHOUPebOUrXlCnGv
b8uQjhQv6WbgHlb6SNizl0sK/ZTE4rZZoqDIR46fMAAIOR9zw3yM7lh+K0ReXmGh
MQ558cQHnDJKrn7fkuG4GYrgECrKMjT+8RJ9mEKUNT+SLjsTshzFisP6L7fhZMIU
5iRMv0dwtbi6L7+2R92YZjdwzIz40GqNWGA57GHkysv8v6CYSrhAw4EN5zZxON8Q
pf3dauOtGQ+Z9Qqm8NWISDBJ0EjX/DXxIrAn5PUym7sl2jDMuzQ+sKEDiBGCgAQK
QhnofajyTzLeOKi3YAFKz5N1NOTn8e9Pj/5AYq+tNON6+TWT5raNpkmhC/4Oe7ls
S89wMV0tHcS9KUzqXxnDL2eUKvFBNmlZAdVptVb84ES94jP4ycoQD0dvleaJwFYd
OQVTNEFJ21eQ0MhqhoL1V0iEbk5jjd1SnFTfeoShNUgZttmnsjdmd5gfJwSb+pqD
37yqa07jniIZ//89keoDNhjsjZBv+oyUACECkGH3ehz36FZqAGRh5d5k0mJhg7f9
3t++SQofjpvuXMhWDdc5+/eUaeA1Oz7HrLq5j5CkF0eiAsTdNSt0NdjwK9+qMOHN
Zf0oFwfveFZc45wmBAYepIdNuq6IPl7jvQbpnHyiHBsVKooPeEPPciAsltxys8BW
mnx47DLLpoUlwK0yBXQnQS6G4YaB3WAIgqueW2sGe/7cRsrsi6qgUgKv3Ue0okkF
nKfh56UaB7TutnqmAvoyVaVi5mw6FbZcw6AWky0j2prsyOSeK9RZWsF/Fb9aHWiB
YLScumywtcxkbAsrjIJgBZKRQbqoLVYh4qtYDh1nDgQgQC8FJiV+fzQh9pq48H3i
0rqxAtAf5ID0bB41ByFK44CUV7LvKMLaWCJAVQtT4HCDtXwCFghHQJ0xA9EkoKAS
Fj+0ZsM/GTQy9ujSyYyvEgE2RN5QeyK8dLsKhqKsMFZQrYdFSidErZjxG2yKwJBr
M8BZohASymCufX+Iogyjze+usxtBYf9qjMxkmCS0+pFCfCD3SI2ovESfm459tkJM
ce8h19PYZipnWo0xrjwYD16VvDxEmSW1ywky2AGwuAHpSpgsq+l+uRo6QFFwK+9D
xBm0Ny/I7F7U84xwP2ft+AKgCd7SK/3vMmvrY3KwsIjJPxUHWIV7VFKBAG9Ig0Ki
sE594F3dLFM8rCeHPVRf6ZJ73OrUVidiG8pTscN3ldC95rLODcPMtnvJDHpKXefW
NVP4LrX0Wg6vYoIlH8wVuDM/D1keU/QbvIQz8Y+p6OeuhNp3VOI/xw0DW7bamAbn
ziLr4CwBHEzNs46dVDe7ElKZK9d8pv/tGwMv9VuOwbxMCpNg21HvUY3xIaqat/FT
JT92Tj9sVkv6VfFINo9BNN7OqQiWTM5HxJEYVy18jvDkJdXosGBa9/iOzKMstit1
CadZxMRX97niApvMhuc1SfZNyccQO0d0sHcqsaB5Y5F1GYdWtrQbdLILCqBWB1UW
uYm8mYzqzBrtbKwrtyXtSOgjo02blQkpOuYZaKc6aFaPcfDvtkCFjJ3u7Mz+5IlP
h8hQeQa+GyRwJ99e7qBXT8iP+DLfXr69/h7pDVO3L8Dd60El0WcHN/96a16+s5Q1
WPQSOp0HZnltZxFZCWAyOPh6Od5x2YHdEXVtUqGR9AQAbT5KHsAL7IPBOeMOT8nV
LwfcMyqFCsI/adQ3Ttwk/TCp3cGrGy0w1ZkpS188nT5h9XwrbhJWi1xst070AAX9
xPIppV2ey5Ygg7fsPXdbEIhJOC+OO/2U49/XIZ8klqW+kVkNO1a8H429o+ExWNGW
pAV6Cx8MfOlql7r0O2tGrOzotOgjywrYSy3IH6uhbbqxxxdANl4pMUq2sM2G6Uhw
uMsmcy4T64aaGrNt/X2/vV0zYkbGHzMg01pHidy7+hT8eav1w/yFAFaCCPhQXd3j
DuKvqQ94TPEwKdJlnwau2IwD21iaB7KTKM63dHRgUvE3qITG8gItRcUDribPN1IW
fuXNv0xExBp5SqVM28cy/73p1WZFU5rrYUJAx3URaBGgWhaRPfvyWP6psSpFi5Iq
OXiQRpiOfeRxhsUcd9kCQtjAaSPvwkYKwac/71XxPZCVHNfpOaJ7GSQ37b/+Y52w
n/WovLFn8OgbyO7NypRToXJIG9M5ii62c8rAt/slapqT/6tHjrnj75Xv1wEoBwcL
B+SlcnLINoi0shvkRMxHHVNhBNBiqrhr4QsbvWnekTipv2YdvW6aSclfbB6uIkf2
Dz/l8lJCTQ5/BSF/te8A5iOxAJwbdiuOZozdWRtknkkKUk4STPJMDtRYWHaWxtTJ
0VHxqlTdScS/q9/SjIpt3LSYYaaAIyxRGuZKq0P0Y1iEzNDao5qKL/QnzE2pllvF
tkn7btkA4A4tplSBniFpUkteNlqMAQA27iPQdkBB1TL7hcoMWvXU2SjcNT2KdKCR
uxx6Sq23b3XaM3o4EXIllXtyb8NfCWomTyBmt35sjrcg0/vuOUC9l2UG74wD9i9q
ZC6JnM6rrRk8ZTVfHeLtlyfhgAH7iYq1wQPAnp+C9D/t+Ia/QrGHTo95GiAvkYie
heqOdWOISsOqJ3a9umQ7LGMxEBC3B1PgwKzUTotOIM5NPQ0uAodGUKIKGUt1CN89
nyLWKMkTOeFJxJi9TfXPDMngWU22aCapIL0lvWDWdtxqLDioNOvaJp4rGpqIsIqn
qQW+hsE3JGO1jpszw0yV56qdRfovzZ03TCeSvA+PB1FxPlwe0xn73QNIxK7nnhS8
J4GHkLJRzlSK38GFQU0zUoDIPgtPyOYvwt3jOnbg/ztP/3BZFyu7dGNkRJR8NVdL
GFEv4GcEtmRm1h0nDMJ7xoa9ZoF28cbb4RWlfNQSmrTokqmq/JUkjqGYpRoLOtLB
nwCJZn/hndk1aHWtEBPcUayl57grWMviOdR2HdLZzAxoF7SgzXn9IXVoSUx4q1zd
eve76zySbdqNk9NLYgeT8if7pm8KqWsvJf4kSddlY8HSqRn78olNm0TF/ko6I/jP
5XPvFgmOBnLfDa0i/t4s6euyhFJwUMBuvbZsm0JcKoT2EamqMO5PcIA8sX4BPr3M
iQOaIJG9W8r/TC4myrvPGCKsW6x7p4MVhHfJnHlUCwyCA2MnH37wv77O4j1xy878
u1xmxC3gneuIQBi/OE0VdC2vLE/mvtXecHaW4Sa0J7a/+bbW0lVLd6PG2ciZSxbk
j5F6N4uKvuMxu1rdNmkROR0KBb73EdWPqZhRhWToW3GlQ+ZUKneaMMRUT7Ufgbga
o/86eQ8uRt/52ZG3MarCJQH1o7JyHaJNAU1EbU8VRdZyHr/lMmz6bdHBBlJ0b8X2
YA0Jzzo4/d35tz+8aoTs4Zvl7Q3znqGR55bBF/elxSXaqwRQWgDfji3kekWRRdAF
t7v0uW3BTURSpJkjTvr8XHBwPLdnSirr+UoiE9XVtCrggVpjizKazCZOGzYKiU9x
HMDP91XuNJJGTLFiNSqaefMcMphiCfccsC+GQjonqboRZ0ppvtd382u4XKlmX/7r
PZ/ssfYSEeWL4a4OSy07kbkqOArWL2CIFRstz6b/w7c9dxA0dZtMtr9RRa/A7Eq/
LD0gZX6kZHV16zr3zFdhtSx4OCMlrKGvREDXpyjk4sKwUwQ/pMZmjJmqyG1X7dSC
b1Kq7DZl9MW5aUe7cTZPqOXnGxlkNZQpi5GWjaawkNvIoTWy0crLTGIGW9kUB+8q
/VHCer1bXl7BpOWU7S26Df95EBqBWosr97EjvJ8wYnr9UCxY8PN7FmN9mtv/1lAo
jRkDLLxcDiz0oQ/U569cN7+QckuDA1Ir5FGtO/ZSzAi+ge+XG3omUZRggEPNGVkD
zIjTrt2EcMAVLUHDOHZdDbmBaSNPap7eaNRkf7WErcVXFaMnIbpq5WC/VIbYMk8m
o+jIhrpkSx/7hCWc26v76UJsftTuVkjhGTX4MZkUfL7gXdahoj54jPl66kZjgDLi
7ipeaeV9Y5lzTxI4nj1JhDh3UA6aMUo6NNKcqkiFgnx8KjhMzbnlJ9aDf92tsRW6
nkO3FFf/ASiSnBIirQxe8Uk2Gid1ihWT/ihoqhDHHnkolpKOh5q70c5OxCxHy89I
PHos2vB5wvmdOMKG5zaEq3EDP5viaEGnUQq7VO1CI2URvAwX2Rq79lZgZXGA2X8F
ZlYyLZZQQezAuZwwNxZqh73TtR0kS6vm6K4cL4ESXPIeFcLFq6Qfl/5g2uzD2rj6
9cLrtCukBmFWLCUQBNinUdkPA2NhhOc5bzA1XTAB8cjtUZ56M5QfBUETlo3DIjw/
487T+GKPhq+2qJiT6e7GOG3aXVpY8HQo0cfounkQh1i4jMC11swg8JMxPeArvQv7
DRMeRTyEHQOynnJj0jjkA3o9Xbla5J4nAyvmRbAm/vxgWjaKxxq3FFLzAihK4JOH
EaGMOIraq+dTF5nUp26PjcQbe5+HfTRl+Y521vy6FP/+/HBnDxpmrzhFRJXW/P4Z
cxsF3edqsXoKzYWqYUudLADSbC5uXlbh94JWkZHzU7cHxfo2jqW/pUk2X1EsMs12
VgccDicCUVJnCxYQShY2rPsDsl3YT6TkzuLkQq3u6EGL5vti6M6Tfs6i5vpJJLKZ
QMNuUtvlG1p6N3GZRX2d2/zrXeCxxb4LsmW2IcrnRtKeV5Ymd+BeGiaavrYOf+Kv
SyPJNaULFOsrjmjyZLnLBS+UrKDmQ+x7vSUm5w5QIeaWdC/7kapQTbXy1C6io2Ul
23qt/FvhI67NOp2fXd/DgwnfIZgD562HR628rZsSpWrtXXon/P3osLcqRYx2nP14
vEEcLjKQ3A2mxNa5VL2iuZGk/YG46W69cVwJWSOmSeP0O92dtL4jxdoZ1aVZXEGg
w4gP7nWiC/wlBh53WD0MUNVU6dMSmW9Z80Pb8RTq+luoCePOVGxLcfVcgcDU5X0o
hZob7dkqTRCFlaZDqC8ism8kycbf+l1SQt+ky0Pchy7PF6VYdbHPgluKHZlRMkMk
II47uBL2xLKUZuFBysoKUpKl2N4QDlKPPQ4zsP9xGrPWAol/igqcl5vI1Mh8raea
QdCzk/NnDjlaWb4pdN1Dz6ATVSOls+XsbjFG1doQ+xoNfXE2ryvfRzMoAVeyPU0d
/tsD+ORkOv3zBRxzan54ABnEdjN8QvrwTA1OphccNeu7UDkXA9H4X6dI90uXXsEQ
mLyeOvJPGkJe/0Nrh9l0z5sta8hgLmDHyJk52LPHoylpyF1tl67nMUKPFI1V4vWG
xJhugbQh2odsmDnZ9SWOli2/MWDZvFozMM1UvUBnK7sMgrLcyrv2NjxcKs78x8F9
YovWNw0EDvpZsr7/4Mnzw+F+MvBYqqvvEq6EF2M33oiCePhmB8eAje4QsZY+SNGd
VNVwPEk6vjo3mURxb2KiJi8YxEc9Xxw7N/0ng5lAwEHJuekq1PtLkDC14rDOBmDN
ZWGYGofi7BdUtyE9VaqCEc6k1nC++XqzvFCJk/0vW7rU0XblfZFUrj9S8frgmjm7
3gEshvLOhBqdnJ5Njho/a/kU1ZGgJ3trL3HBFlOeRwCQgc+k108Hx3Fv07nFc9cb
xcPBogVfjluj8uBnNvx0GJzuW9rRRy+iVIsU3f7eb+/Ho9ZtEk63W3fcN0fhnkbC
109LbvNhi0Ud1ZmS2VFbeqC2hg+IsxY4AKJkGRN+K1Vf/WO3S13PkDrXatjFLgTV
AIl2xmFAkYW9dUkmUGWFDAwSIfBydno/Wv15PBLWoBNNIKjheUrRNo3B/kmx6P39
h7BL67ZuaZ5LHP2/AJhyeoYWIeoZOXR4n3j24QSQab7ldlgT1YGiUffhj8kFCxqg
j7NcH5YkxyX2Nu/jctc0czdivNbWVvK3Kp17+pUccuOv1i39dd/XlMuttGH8uLMt
P3w5BmX17Cbg1l3h7AgX6/fI0XJ+Y3qJgjJha+/6nsfTo6HlN0eS+wO2EkR88vF8
3tpdGZjoNEQ1yBjxO0iqn3h808ckevJtIHGy++sDn+3uF3LNuDwkG8Fp8MNgvAR0
GsrMdOYVv3NbjQ2Cs3j9vALvqBqZQqp0pE+suxlSQ96R8JUb7uPeKEhXhfXQr6np
a1BHcpUOhOgJZ+KprM+UM+B3cNWHrJc5v8D6NDP1sdEJUeS6aZa+8xemZonLqtT/
Nj9JJJqdBx53gRcYzif0eURD/2dEImot9xIv/QkGVE5qf8oeACdFpChbl//xOHUR
kNHLc6Oa8sMxgjih5+YYYw03dpcXQystvSjAXv2kWj28jrGZAt+fJlPE8chMK75f
L5JEmiDoxXIwvtduQQjOPdjjd6o0T2fXnLm33S+YgqcdUUJhNVHuBn761xRHkWK3
CNdaY8e0+luzBfLLGSpudcqyCIjopMR+8eaGd3US5OXOPjFYFJXIIQgrY7LNMUm7
4oVqO88gLPXg6hfYbcj9OOUlGaGU3ocEkcmxjuAfGXkXzj9NgGvJOXv2+vqu03k5
7GWeOymGiNMk3UH4dRdDiuyjZzBSZGsYwR+J4Q/xKEV0Az+YR/qvBEPuHnCUAdbf
p6u7GzUGQn4y0Fdo2UVgdc9J3yW7d9p+vcQ3X0ItLxfNABrO2z3yeVIcT3BZPobI
zebFQdw4ua95atkdP/SbTgUv9dakmh723UW/Ntu7zw05PNvBXQmWaWPQMCxjDDQd
fjDqzCAzF0JM1P9tAz+pOdkYWO98FGUE89APeHKtzcC3jVDjOnlSbdn4ecvclwH9
e3afAjzrnfjAYsKPbl98p7CeFwtkVTfrqAMFipocjjPzsYC2sL82dw/WuFmz0vx3
lRc7kk49h/U2c9fjfK/B+nZ7DykXOyY49DDvPRkuWkSt0iEwr7h7nBjouNSAd3ps
1YxbbZgb08YqXLDGKuwC/QN47AGIw5P3JclhMTikwZVXNagedDEuMEyot7G8mktW
VR6NUsQ0IGPIDFy+KaChDrcF3MYgIIkaP/wYO3s2zPM42z8OhHX6Cpo7WQJgu3rX
6D4h6/n/kjcB+ZJvRRMW+3oAujfr47CC47zN4AeDBtvmg1+CC3hb3Ld8mdYDTH6F
+IbU+18a/yg7SU+370keBeaj9R0pAHCec8MogNRHtE/DrwkmIX1B5gXX+MMD/jY4
J8i9DlcYi5vfMoLyqMCMoBwqniwS5kdQ5jPBy5z7O13CnAsV4JUCPpmLl6NJKH+8
LlfbJlGkIu6O0NiPcqtS0M4oZPXqLN234+TZcLLg2utSXg6V2NMSLFHKpVEZHnOw
vGcIxhJVOJdDodV1MJzcYOtHQxTY4GtwHC4hLBXRwd9M1xJtB0WyA2ID+1459D9W
6ajJnJnUkmf2x18n3kkY5UkBEhXQmeuqoNXL17NzqePO6dY8lT9R6kigA1oxRnYj
cTGCf+Rk64ETJLI18e7umNMKsaRuIFCR1Ey11Qv1cZLYbNNOawHnsdrLjFB7/Be7
qzV9mqULLp8ZZ5rT9RuwYbFVoVtEhybKiR43Jh+7vyDZo690fjbTnUnmCbZHZC0v
lgrRkiQ0+hCDlumlJFlQWAfBPaWZYpYnDQuQPZeeafgE6Kr6JI/rrczhe8AjkQ1s
wrfSDTKfLWFfOj2XxNU41kkeS9e3OQOGbq8E1fbhmryGO21EHq+g1Lqcg2dMukEF
s6CerdI46FUnDizTswRvnVr4HW433w779L3eD4PW0myf441dc2PMswSpUgSpMLHd
3U9PxJSn1jOfc1vLu0kOJ7T1zz3uxf1C7saxB0HXashEcO+KcZBb7P6lHfcf/mRX
e8vQPA8qJp9rmgO7zKJlgngAfYzt4/SJBg4VPRCW0blxSjOFrsOJgjI/QMGOheho
fw8R5VlEJXD8Z+NyqdKL63+Y5dAT9pO53dy1iV/QZb9h4tIHw4LhvW50PyfCq94P
7suP2yBw1BfWIio81uqXhQGTPhcKTIAiFZcUeiKz/MOjY7gjN3F6wlCP80E6q97d
xCGsfXkHy+53drSY0AoNwfE4A/imfY3829swr9KLPwNlF+IJXsVNuF6T+dQPbp0W
f/HQQfOoGT/CL/YTnnK+pPKevd/tKm8rNpjng/UtPLeifz+vSOI/rq5aKRTPe1gv
wKKPENRv5406L9HGaByojmXhPwcwSGEZM7niqOLgs6X2O6hSSLMuo2HFOCEsiZXG
Wls4kwHfe5KF2CrvGIJutij9Z3l/0L0PjGMj3FIToEZSit8q6SBudGtCHiFyyXPN
OdeWindNUJEXXxQswwQgve1xKQZKAgDePS7803fQvOcGa+85Bmh7dH7DG9zJHSfA
Yx4O01wQg1Uz6HiOUmlnhNCo1Bqx7b275WjOfWg8wNLrBgySA+WhfX5VfVJOa4eR
n5VnKfQ6JZLw91BYRHKheKEBZTZZOJrGaa4H09IGxNqp52Ca8qMoUdrWnB5SHD6g
afmzedy6m3nTd+syUtCuovNdhoLSrHe7TdpArcErAtpa9GYzfi8bqxYDC5d1FKgr
x4d2p3EFfSZznfS2LTZbtvKQIFiAYjLgm9aw75MZLa9bzp1JeOyxJX9oCsjEgRiC
bm3oIZ/EW9tlp2wJxp4hCEsubDqV4Rg8naC8E1J2JdXrI+2ckS7wQNrT09f1JSPL
WCE+Ni9fxdutWd2WpVUeeGWWQRLP+2Ilse3CgzkUDsbYqW/XBKbFup1D0txIuD0I
fZqA9Z4GLF86QZsh+uBsTVEpJYUm3QNSn+oAQ0pTQ7EKFQGojn9UeoLJABDQAxhA
2Nct/NsDiO3szOFM+5f9y0DJ0tIHa1bWSQiPFICxYO4dP7E325J6YitsAgM8rEtB
OElmc0EfHFDpbTTecI7Ye3T6Z/2tG3n4HEHpcbbUiAJfRs/+YCHJEzp7VEVNzwd1
6Vjh0Yr4f67/X1YzUjKMO1NXoztewyAPWbdggVv1BRPsjR9TP77ItYFjruqrH1KP
M5Da3z9xKfOJvfPsasOC0P44xmmrd/6RoQX9SQycSBhu82fadaW8IT1hngPdxb1J
sIu6eH1gWlnwBpZWyYADEU7AAE16BFlWB+OcWXIqmgp9Xon+XfF19t7hoh370Q8x
IfSL/9xxchgEqAgqpqVoX0r3onpTC3MKOGqt+rmJVClX13++AFwh9zjwVhsNFI1X
kA+g3A84gqLCGXkmMJxVbqJ5yRAXahYoPff9OCaBWkWi8U3gauCJ9IrBZdE/vYvX
FgEKwxbEtEXgfz+UX0sGT2ooDu3sjP5bjrCfdS+kaexRKsK2L+h9ARM2zvQ3vW7q
YgW4H0d5oNaNMEXScngR/LbOhyZe6fcFzXfBlE2Q4mKsf8KCVKfLyJTP2MjvbX5n
ahSug4F/ShBMTkWXOrgD5ZzIsvc+k0htL/8qoREc0YfG4WTsSTh+Nyqc6z77UOo4
qxdMic8zr41967ch4KwphLWOwwIZgDQhYtz2TA8TuBGTQZ/JN9Tvuifur8tGAS8y
QMpYx3qM71JVyjr3V1YF8ThFs+SekgDJQhKu3vGEUzsXN3IKrYhmVV3b8jcxgy94
YHK3UmQXSW8jZ88fp2r/KkqVryiYLxpb9aoEl9/1nZhdWXyhk7i+F6jjakjrHBoI
bWBdTXtQDEFFEJ8x1x+mpWCSAm1mXT0ObWcxF6cdJqZNsxh4wW4fw/ro37EjZbjV
GsZ5uEv3lNhknCB9T9ydbV7saUXGlIJPQLx9APCY1iVDmhrcyQMzbYfQveGbCRTg
8kq+/OPSYkfZc8NMX9VRSGSeuML9fE/jBm2rIAgHb8h0HgDV0gAMX7P1zNbQbm3M
qRUBgyh5RBNFFtlzYYcUk6dreybuJFCsacrPDFxvPF+OJNwRASIrwZinarsm5Slw
PNriP2iEksYxYwNe1k/iwINEm+6q6mJ/Ffz31o2fE+8R/bJ94UBBajfffoUcQhkb
5sVnLVpPsF70jbUwygZ/C+1PhVdpqP6QQ/fLToqIwcf9XQUONiOfsRgUhtj78qp6
uPID1yRNVtUZPgIGbsa6i5lbxDDCGoWKnyqpuGhtY0O6DBivayM2yQPgLrnOL/hI
r/NtyO2Q19fqrgdykhYQFVHRtkNE1LJNVU4oApAbvFV8EjNakc3K8Gh0l41rzSSo
HSoxjyKt+5CbPem7nfCNI1qkm1R5s4+3gCoWpPR5/ZQ3Pwoc6FY4togf4tPf0d4q
Pe00b0zTwTWvMVjDaEnybU7axK3oAthjUI1Ie7FLMV0Z0wyHD4CzVPkmzHJby/Ii
JMNzScyJVAen2X5RIVFY0aPDmEvSQk+rJTocYZ66yUuRwnd8CtOp+ZDJ7+MhOY3S
4CCcLpKCH7scdvTRaLlMHrAgsrlJokgDpS4/7hzzLuP5S1rcyfnYgw0m3Ud8XyOE
t5YjhASD5W22WAzfg01eN/I85ptwITvKyree/F9RpsEhrUJbLAEbhCr9y9SvUPJX
QgJWykJv2MHIXiZJSrQJPG8Alcu8dj640lMAvMzxKIszMZdaj1+vJzBqGH7XxEa3
NL8t4kuRhgRFEj34sd+swc2fV7ksfK/9gcTrNmKgqTyX9iT+jJHbRvX3K+XwaFHg
wVLPFlbpywvJuN+k139o7M0z4KLYv3LuenHcYN+L4d6YT2viPjrl9KYQXlyevphO
X80NSbRmqO8oSe6Ml/9wlQCcA2Us1Sx4bvp+TFaDzx04ThGwWX742ComlxlF/EZx
HuJam3OGLS+QQ85APhY/IlzC4ybctflAuhuUglmiZiJL1jVnTavDMYAHqqIRLspb
9qykIyFpnm6N4mTx5GS3sJFRimVXDh/NnpL2w4Qa8q1voqwTSeJaQzifbj55yc4I
LL9ojJwU25szv0FxYMzIAFWoI/djqFLlp6O7JBtcv9a11xMFzbuY4ZVFUzAibrSG
BXV7NOsUHxn2tbuvzZSkD44998+MvFQrQTSyasL7GJKG0+/8CqvcY4bM5ZESTiBS
yFjIOIspa8BPRestKf+Yh96HPg2FyI4nYmqNEe19iizhCJIcCk9DP3qX7qxG6EN4
JjF2OooVY5c6r7BRYZ8a2bsavHEK12a9WcDRcaTxgtFSacI1vPZcatiVHZwYLFru
n2WijKkgoZxDHywsGZGY4h4rlvhq3Q2/wJY12VdPEAlqkRy/dQWS1uxDV7T3NB22
sGv0ftIW51pwWuwUaqgyq23MhXc1ccxpKMNJhw9+XhNo15BatsiRQrTOrSviWJVX
Se591dI1M3mA6TbCuldoj4GdsSlNxnsGdU9+9XwPqrKt/lKfdNuL3guodtmIVwMx
OeslZ3N5JHDUrzRmvnufanGI2U2Atn6sMkd+hAKWhtue75cH1TF85GXUPe+7hJGC
ABMObUDj7Lb4GA0A+9WbnPssPVFR2BuEBSh7nG85wLUihxRE+lQ7Ayp26UTbIHfL
MJkbi6drim9ytN3/qmO6op/0P3bbKgIRHbNgPR6e/mAm9NlyrXdIzhj0LCmdHwPQ
cKj9Yvkm5Hr02cmNbdRENLdOo5iiXA89KC+btaKlkjUnPVGsUB7gIUnpYrFOhG90
5W6VgQM9FtqQ2Yf1YxujKqPjU4GjMnVQm6UQ9cVL+ShpyeT7kUw+30I7RXphMQ7z
vFQ4ZAlOITL/pm+znOIgk8wNTDrbzMEbg4fyDQ9YCATMZjEnFUpRlv8vP9FwSVv3
d8Lp49wwHdXH2QboerehdpeKcxygwP2T903oIs+6kJ51cxFgL+NHdHuO8BoZ3QcV
TcEnoCwyg6UCd9l/45iyn0f20XcJrk6brKsAFc0c/VXtYDYK551+W3AAmMa/uW4p
jeT8uYnV9AmNbr7tmAX71cQG2M7V0NoawIA0B7oIQwWC7wc5e3vWdtVvEp+LRg6G
uzJq7ArlQJg5tkmaUVDD835Cd25G9fVJCBWV0BSaLxiLbCKcwNwxVPCWBV5lANF6
kfRSnnbCt8hQwTFRCTTdSdJ4ObgWXKmtVyB7PfuRRSaPhIcW/ul4Twhy47zx9k2u
lCG5sJUFWGV/p0w9gUkzS3GWKYq5qTcZ2NergJGe+9pRpzCO33b1EBNDY/V6HreM
sdMNpqqeKwZKiE3PlAP7p738TgspRx9XEvzUrlvAV7TLBQvJmc1nx9Oxzv93pzmM
dAF40DQeWMeBPr3pX+uAU98jt1G8The+yRx0tFnvgn8otwy3pvNLesFSWnZh1Bp/
6v1rHoejbHLZhJcG4dOBHrvIUGqkAHUZigMT8LjfDQYgcZDz5J0a2d53xxsFsRbv
BsbdY1MGLk5QojoB+SqIO1ZhEeqPnuKnoI//jEyqELbxOAIrlgVk1gULmqNbv7K8
zHIigWX7+oRbIidEbR7h4WeGk8ZWud1LcC8edAQM53GtW6Y6V52kPrsMcdjUQMjL
kuGy5cA9AuYNX193m7/9grX7hQwwVP9hQMSGl31or5sVVrV0Z4r8UrpC4O7hOVaJ
NgwJ+sSqJTBpUvGnwGF+VNswIzfz29Vzg8K2rweu4Mge0LdnYA/TuugZuFijmiOA
f8MJwIkFZPwJDSjqFechJfiKzQISz5tlX0rydsQLv53T2jddGlaVxH3rCZCdhdcy
wFpN8obSJ/WMA9SkzQCou5eIQ3FuEO3VdKec5ZyQPvEqqIKwlNfKXHgllC7W/MFc
IRSmi9KF3MK/0tnwSl8GtMIkvpU0RnRYHStwPDxMrtLBgozKOCzNR9lNi67IcHtD
+Jtr5UWP2+3e7oLdnkt0Q/wqjQMjDe2HRrCbUMvhpqHusIPZr6khXFwSewyPYP5X
b1iIzQMqV0PQocm1kwIKY7DjTHo1OrG34uQJo3tlMax70BZIPXfvFlLEaLmoHvZQ
6eMaG/Oc4StdzKETFt5IVouaEBDjJVRoKX6zJAAyZo1/rhQZqoIEZRSJd/6yeFLI
/mqK+T5z1yhoRVBIr/v09Ptr+mN7ALwUWMH65RX3piaNodx1J1jAzZ935BOvxUxu
LdyA2t0B7utYBp6Odkwv9TIsGFwkr1gt6lvzxeRImLL/BNtWWBGW312mPpOIR9oW
lQEP5ddyp/q5/18yuq2M67ycGYi72SeiY0QwdX1UYmGueBQuxhOTmq9Q8TPMMVKl
WTCcfHKMKFVpkqDROFpCgqHLn3r+DZ6AdoTeM+u9MohYCA9YePF4m6/Qo2TB01Fm
AHGzax7/keO/NdP2qUJGP2bVZ68jp8xYTboY/3Vxdx7yLzrJM09cVRruzMPGDxpY
OaYUDC7Quk3wS4JZT/c/BCatE3W4fYdH/WGcDCuV+Yy9HmLLKxPnu9yajzHzh+wr
MaDFfSMh5wuI9Bftsfa8jY8x/rwr/uKzuFOpkJssk32mFtJ3hd1BxyJ43vCwOsiu
5slrPu/+t81ptRHSMYHDU7ESei/vH1hr+NqnbDHBWoCGBdneW187Q8vSTXQN7mqu
zRyWxBogTubOV/3C6t/tDKpNFaZTXOiY8T/jtEgaRiaLDGBQ374W5DJ9d9qQAxTr
AozM9/jLnFg3itwo2wOS8MADdk0FcvXeR0zN+Cy3APxGe5ORtURL4vFpBxjVXvi4
4zVQcZYhnCHCqqqsH8hl6XngeFKnLzOA81xkl3uWEUto/haN1JQ/Lm8gmnV7k9Mo
zgqninR/Y1mR4zEd10kfe1jTy3rPhOmmFpGK9ZF0LvGgUf8JnB2yh8TkKZ0WhwPD
q4VG6lOyvgLNHg3gEILRU59axSoKuVzh/A86hyZZ/kV98bYe9x1ecsOl+9XK/EhT
24hC1M/Lrvs3Dc14G5Swb3e488048wLpkvIphI/zUMlwjLjD+p2TGhdbV+1FSFao
q4WQKV/fjSNMfBN51cL28ymNNMerJ6ykaTiBV6ipg4JBxbI6akTAve1dhADFnzP1
SiUAGBGuUpLNwU97PkgkIfIfJ29rerCjrxVQDqAumQBoCBDV5LycdCnU7GiPTOir
vyGcU0kH7d5nYYEXff+GaIMaCKTutmw8YplTbLURZaW5XY8J1NFJ7975ljR+bkSM
xhOGC/TWka54I5h5XPYbKDt445eB1tE6K8c5mvKZm7IE/fJ+Hr8sU6cps8pMKjE8
Gh8gpkYifzKW8JNNKm4vyuPSth1VZMSdZYdqSvW5nFoigymE19JDhLc6YqYX4rj+
+knOzKMuJAegUC8Lu04rLsBgt0RBYp5vYhyFYaKngh1u5EcPn1Z2AKSDFmpPOVT0
qjSFmxR/xdl1ULnva/Fx02QCbLZCS4aWc9Uy9m7QpBtZLLxlf5QfmVvlVPjseuuh
XnFvAC4tOMVRgI3j5Z0iPVI5bzvUMI8qEpCA4n2cTj2F9LZVNsEtPPUJMTTF53Di
HtCKUlgyZf3iFcKaFOyfsrn0fh9BPZtBFD8zsoDwXZoPQ6JlAZCk6PtNS4ISaDFS
P220IC7pYSunieJZRWpEngryFagMl6P8XpcqK66VcJE4yCmmKlvESZl8S6qX1yzn
Xk7N90Kkc5xMDgRjf5Fi3G7vgAxD5s8y3HcJqpYw5zbSX1Jqno5F8bjNOnURBoEj
oeQw1Xb+O3BpcD2etvUx79PZlTDgHEMXyA71ScdTGCX9UtYfaE7BZek93F4GIFo9
n/CBlJT+W0DYVtE1VM15h6LJdqXRFvVc5bhOhG749SIU37FNt4TUmdpuPcZs/hyb
iATH3uAlDpHJaf/cSkE33j2BwRdsPMUCv0nc9hT/FKOGP9C2WKyeJB7Mc1WpWLvA
uKbxT0DdXDRBwKlmH29rMma7RcZx1oU2FuamDFuUWrKUiz14lT1qIG+0gOxFaqDc
E6Px3cyDfCCr29ZaySKK13cs8sHHP6xu7ZwFVK4IET5Fci4N5LvEcFueeIopXYJN
UmWVI0JPr11K+qgYSTaGPqomiLT3wMUAYCZvFYaXPjhwusQ71mcF4b06DcFR9Nf4
eJCVCfD0svFanwLbzBTVaP2hzcpbybaSnWQdjuKiRycrJFKIowAyjfTBhq5ipY4B
fO/Pevo+1P05csJNerBi7s6Eb15VBrEvpMeih4CPOY8RrteIfulH+f36GC5nmI0O
0omk88l+WxeSjnM7mltI/KZAwVK/I8kw2oC9JtGgz19c/pko9CwOUrg5mF3ToIT5
UjuLqExa5acPOGGX3TmlddyN9rnGeothZ2gWzOjZRB8AvSqtV2tYHEzzZPkIBzXd
XrgcyuVb01nMAA0pD3w18tBSeWdELy7fW7q6H18acR/Vn988x0DUZa1BqAcllvWP
3WqBlP7t42gen0h7Sa9Mmb8+Fvrk1IgP4pjRjL6aYQaPWJneoG35N+y3ju6p9Fiw
Iu3KNZXPw5+KlU78cG2hl780rmywQUJG3Z/Ic5FvTqo9ptf48s3D4fCVM4QR6nj5
SBymiP5v/iPG5aKPunDorkg3yau8plkXg4BdQNAIupu1xeYL9OgBZg6zwOP7KRtb
Pdw6u9bDpxt/hxvFDDnLqaXRdcr12VxL4D8vL/m5vEB9sHhsaR5YWxu00dsqimgB
zTl65ETAs/rMS8L/96bTauDgLEWwWxx4R2V/0XSO7LJIDmSv5Bxc3Hjb+5k6X87I
F46z2vavT2zujJYxlYIcOi3K5HiI82gQPnHAZ4/5WeQGAUPuwElqVDMnIc59jWG9
W943YGbFZHaMRjVRr7sTsxjNoynP/r7vHHIss3izaz81CvIhvmXjblkGNnuo7fMK
WDOh7T/NlT5t/+qlqPTKGbKie3c02ffYbh4ZLCeJvOAM0FU9ujUd0d1JgXaQpV0y
N2oZneIDcUgkXyZB6Ao45tDt8oA1u5TVyv6pEuMXDpnL4fC7SgYrkKolSe+goSUU
rH8FMiktnd8ficzum4T+FEDwFsGVocq9hx6ZOS+Ik9KaBO8AHhQR7czGokLRHpLl
Jqs62nHosjKY3Zws2H7LKrX5Dm/aw7zRmnc+g+OdhgcNC9u3DBUW7FH+5IOiWDK8
l605cwszYO3mWH2OBCSdavPcrcnm68ltZ+/VFl1JYhrkuRjJVYz2g8RhDyetS7kU
h3VTNkbU37ctx7qAURx94BhT81HTwfG+m9Ov8wLJUDh6/pVC+Zzf99nb0q1GU47b
PQHg1NOV0F4+TnG1UpmzrcrscVKyWwceTV8VTtdLjElBWb4OzGvb/s29fnxG/8KS
QJ3CszXEc4yCj3hTsLC8o8B7uizMbCU1ODPWC4HjntHwMMfpq2jEzyKYkZwRJqhl
0Vf4RFf6mL28HUZEwyqPYblBYA9WqxLkc09sWaESU/c6p7HOtquazec4IfeqVHfw
BGnImGhfNaZoyFEbA0LP0frZg6phOnS7Fjy7icx/PjL58v6fCyBaafvI7j2U9Arv
J5iyUEWYve+aw6ttxyL5hxtmygSQp9lcoORPkY+Db9JSrarKg1+8tRBbrU+JmwnY
mAU7EN03HCNiG6RGIltYkWh0N8N159KVE8UP/+qhfo8WRNAA5RrFGwCqKUpL2eff
GTkPFFAsbO8tY3z4zMq7NHFwaqyGirHERzErzJFIDeT6cenacttI4RjDT/euzfir
GbeyzflxQR9NH2sxFs7e2h+nhp03agHIphqMDx4CMka3V9n9fzANoaRhmJbvRIxb
2fk0WauR3N8BDOD+7CIpnYBGfrF5t3n1eppDf2AQkymEWiohl+au9jebf176tv1g
792JXZ5VbpLu1HDcjh3Z859adwuNM6KKKvIfDr3W2O6/DSp2AOV7+y/O+VuNc/L3
QsfU1TePikRPNo6aq+w5RYCMJvUGb6JrOcAFZ/cgRqDcsfpDkgGwDFn+bTM6zYEy
2nYZTpDTPyvd4ekvKw5TX3scdTMugtx4Amlrm5dHpIs2JK9u7U8Fa1S3PN1xcuS7
xmvsnawZ9tDtLQh2FY9MMmCoL4LvmDng1qmkJWInRG3tmr70y46D2eZU8d9RSY1d
PmG6JiWMV7toMY6iekMY4fW+MB0N9c8dCyy7cACmCPWm9QqvmeMsAsMEabrW354p
W4o0EbGr67+wqV13NS5gxClaIyPX2DwqfwPl1tr+dhXBBOXVw4L/nLLXRbhZRJkt
JRPobeYdJeaTV22UeUl+a2nh4BSMqeHbN5jnOzKFLPBn9wMKXxy2Jc2ihlDbtMrE
CRt7X1BGMOgrC6Mt5HDz02rb8qWcgHw3NnIRQIQe2B3f+JAXllDS7AStHt+I2ETX
t5LnAL0X3jIoGki2B0yhy8uSyGKcCAauUFajPOQHlJxfNfbx22n63njP4GSlGgoZ
GvQgwPpuAyzx7xhRKKcXfOK8O0KOFjIEFv/ORiFJCDz6znb3EBbpFkx7bS+IbAeV
pYZ0+nuaxadoYfExQ5HScLOudOYnGsRY0UsLVTsGLqbUrlaRyFGhZMAG4ctKU72T
nPTCA7OeGAGEMWCKm0CQzBoXBke+MVGpj3QkUkI7rdv1RUcgVQXozoekdTlTcBqL
2Epnomj/+oZov0ZncTB3hMazGhfZcG82FOFNJFwhogZeix2Rvk75aycsrpoQygeb
t7zvdcknCse38VXY18URprYNE2RXFu7ThWa4xTVHt3akLfAW/eGI85NEeLWijHe0
7ciEQ4/TiO64Vfz/wxo/pXHl7QND5zDmHMaP2K1rGURuyAZT7G5vKouavPzPVfhJ
GJPI55z7v5IAHDRAgMv2U2Je7jx8CafzAq5mmFCQioV2yM/2j41O3sPHurweafyP
W8mMma8rDXdIutkA5j69/0+bQn2qoqQQhSsv01FLDj5ezNcqkmkcdohJrTxa8a4l
k+l7ViEuBWPzv3e8gdS91X9OdjEIKS6jmq4u3Gp7VDNrpO/LMnxofTuUHpcnUJjb
YFD16ScabnvtKjBt3xZd8FEzl7OsaddI7xYtXyjsRibovbe4hO0wvY6zfld+d76j
ABSJJzHvxbqaj6NDRnHTL/kVhm6KR8fxu85nOzc6ESbLf1YCaPs0WKSY3uTw32FF
8gU6n038q9YV6O5CcVUygaquJ9Y/+ZdYD7OHMzQCFDbr7baRwAI9rtCtLXX1aI+k
mYBKN4ngVbM5XH3FkY8Ni53fv2jMlqOGTbtPdo/lPfzw/xXWUTEUxPW13vZWk3m/
0KFy8Xr+/dP6LJwqdT87z+BxBdXYKY6Vg6dpfRN3WH/80/HolVl1SVHMMvPHGY6D
JjJmx33arHOrcHvRTXClPOb8lIzg1qt714+CgZfAOp31pjBGOSP3xaSUZV0KpXZK
U+nk5dFqqODoLvfVojJmGbB0RIkvTkMZ9PztKHfaqRm21WwZZc6kdunv4qAjJXy6
hbLK+ruN/H7nAtomVl6QPVKL1a3gkgFjSkBaU4F3rTcURj+JGk7aEhLJUwckVGpv
3H0BYKjOujVQ5Ug+KqQklrKsip+uo577ZgBSY/WCZfJfqGwTeG+zcaLS8IYdnjuU
sKsC+ODvFypI25Q1kisPdf2dF97Sbuf97mBTxlwoo8vmx0wxalJSVSEtIQpCvnnL
0YCC1Vq3UJE+99s0ThQdQBXvDEEwJfmuQqcIoaxEQqzzcSO6wDWxnYvby7rpa5VY
kU/UHN6hSnYYf2XnCEEYj7WtqtJeqxNbTtmYEJUiXUIS+yUSF425tPK305V74lj5
0D37ylYYlvea+c/bl6SN1SQ0HilqfS2pFwI/EuNv8ATipez6e4GXeoijWlsokCOr
0CqTaidalqHwp1ng9RJnkAKTOumXyxiJGHI7nnILxpgyQ4r9oOWfcPefYkVXaDE/
yYREJNibQD9SmBtOK2K5eF/r0/933aWnwyX54Jp81sJ6IU1McVGAJl6KLKJrUcXU
DnvdENfzto5KyAgi5w0xQvQY29+IYU29qlXa5MSAxQhB2xFea/23eSLl1K9FleRE
UToGQKIV41BXz/nxJ2Re3XvE3gWUZNFMAhq7s76cOwffkytYiv1m2I8CEXLfREdm
4OVPmToHYa3SoyrMYJD7D0HVul6wtWABu25madFSTYlQ7poz7n5bT4jcgU57kUXP
OfVHEcxohB2ojEkV/qOjijr7G4Chp/KXTCplRwTG/W6GDnWllPcjBdHc+AjR/KIG
6B1z0H7ETFrqVRMYWlbpIJgWDjfHu2pGXFBSnxJVt402KRkKrMkMhT1k/V7U02DE
j3ZgxETgrG6kay9OsfCO/k1YbyKMepBjQpR27i9BbIBS3sJy6fpA0NTJaD1y0vZO
yM9mUX0JLuKTGXOi2oHx3gJvpgJb/XjMkGN9IjXSj1AArA6zKrHkSiZUnaaHDO6k
zymwbLP8A3ktgw197my8iYvLOlyefydIxOabbVhrR+cCldp5bD/t7U2NATh06cDk
9h/zF5tL6prkUD4o9v0kH4kw0MC8LRSdkPXPauNlx4OQ90LonqiTGuwvBzEC7LGj
2hT2AnxHPE3xK/wvkGApasvgfuTg9euZqLmbq4A3Px531lqOcc0uW/BYDO5ZOPvJ
+WkSXYnNbuhlT3IIMFI1VcY/MgfDUGzS8Df6eX7ZkYGF8JXpNS0ohW5jrVWM9SMh
0o7pCZ5bYWyIA8XU7TLtYxIP3QSu8q1e7CTkxdHQIYHbOoFZCknXosZ66BRNdfST
zWsZjKunez5qEYnceTwqBegO/G2lORoOlhntHuFVgP7vfKhMf/gtlzZlNWnbv97E
spg+xuML7XmPCM/YSuXgjmrhW8tMMyOK3E5Kh713I9D+mBLK/IS84usCfoQ4xrVK
fNgGaHkSUW3n49xgLjR7uhHgIQFLCGlWnPC4zMTF/q8CAfHn6PruWLSxxTBTHIa5
ozRNYm7HyjxUQGwoWw2jnjAwiACf9GHJMfmKP5Aq1rQJC0Yh/S4WSmbj0rWPmhpU
P+NhSoEEh6B31DoTUhmS3CS+PqP87Xr/qEoo+/GnJpQ4RfowGnbs6asiDS2jRx/U
9ri0+PZ5F3Br5V7ltSvzGC56WXjXr/THKyq1jbxrWoU8gEOTfCpKQgaAKGdvXpg1
DCmpoDsujBjCkoaSYiGmG7sIxkafxisqjEuJDw5ND3rf9saKOB+tTqRhKlarM/8d
tD69HmNTwPsKr2ISMrDqXma+6gdSu8lgMNuym7+DTRk7AZtCDhkeodHXiSrCdcxN
Ie5tPTwJVcTIhsDR6900hGfuGaJBynCaTQwPheDfQxpFfGDtsK+Z9gr2ZricN7T0
V+DaWQ/cntyVTxKaafdXDEa85KcOcQE+lgIqKvqUv0uvpADxkNPg5RmN4Fr67tbQ
nt8v+kPSB0xYSPW0UOgUv1WAEa+G13ZEODsPxF1g1zUn36jsIXQYhlvdHdXCLZvT
5FiNZrHNoLKA9oDx6eQO9tfaFrc2o8CEkuu2dat68hkuZvzUdXGkwzSGiz8NyHws
1tTp7qNdobBHxJ9jCeh+UBntW0w6W+wngAc0zFPc5xIPGQv37UJr6bOpJo0+JiCd
sM6GyCLUTSDKFpl+U2m7RdUr4RA47c52vnix2Ys2xF2D4HRlk3Z0MT7qknryaSbc
Ptj3GbYQJ8Vl4YbtTY9PuoboWRLOfIssLUa2nviX8S2J5ug8TererhrP7pIlKr3f
y9Q4KWQOnaEGZFVPW9mB7zM+dssb5/S4E+m6spaV2n/oPlAysHuGsjkxvvRHHsBx
A3g1SgSztkMtkTOMzcN75gjLUB8+jqJnVgz9wx22Jw67H6bG5O4tKeiICtgY75dH
yv9EEued62d98KUcqYBw0TePlT78CNnfu4FTtYtIdYGgjzkTb07MxNwWmbGuPWcS
3gzsUbOTwy4mkcjB08EqYhxI3wNyq2QDG5SfZkl1wbf1LZOofgKym7l73Pnfhr8j
2rf1uE0gbp0gIR7XX/S/PXgpdKzHR4oskZs36A7dimlDyxR7dl4dvFAu7r7jT1cB
iZTP20BP/VtbdrX41sZY0hXUwkMgBdslnUdvg2A35+aze6ywJWVxMkOQD3fJWk2L
Nt8mGt9DWTd3GXgUNUCW0eulz60IQJ0SbKyvan3dcRwjCTfALdyTj1i5EyaxjIEe
7LtNHHqtsrMQulBXjcDKceFgfNH2UiiPYYwa1HrN3a5LbrDQTj+3boShB+xlSxSR
vuy+UzEiqna+tPHd1r5gTNaQSEH7zNhkd0CO0Aq/PNlrSWLbBKuiYA9Wwff6v7ps
jwnVtQUJIsGZn8d7WnpWZznUWbQDRBcs3CB5xPhfBJ6xEwjuAMw1fJY8zIHzUUnV
Qt+vHFQ3s0iSyCVjypj+yu39G1pb6gtT3hMnr3QpOi1zSE4E4MPlQnRmgtADCO/4
PG6r1n7+QUzkna3byjBRtK1OiMejIdiLgTrm3EOnXzy6G7frhTPVgUuOEDIg9mq+
7PJKQUnrGavGGjcoKlx9b60X63mv7ZbkG74RqUyFmhL2qudgvr8ouIUfT+CtTmwd
mfcVoBGxdys5Yx0j+NT5YaBoT1xRBZDyzEq814tv5FDYBL24FJBgNW2oUUYZugtJ
wXZYXhoijxXk19JEFf375OTkzY76AL38icIZzTeuYU4co+gOmsfL3LztdEAVF8DY
+2LaDdDxXWV4EbWepxjmNYFClr6ZJh5WLZNDynmWZYR5c1pDVR65Op6K5VimH+KR
Bz8+LdzbACEku0fqxl15H1PouXQU/4G0Xm5nqrqd3taF3IwLZCmIdNMiE6CUlqWY
EABvEGLEp4CFIYdN4k7fidlT7OjJaDSQj5R4S07IQbEpVXzbSaAPiILXQfvK4tF3
hPHaRhtPfsxg2vgz9YsL75ly0TzNPZ6tcVs1HH0Z8Yo70Z++k6cD0yr2fv3YFcon
r0SbammNn8CAdXDyj9EwMIL8EmpXoBeGlW+EEziXssHNOoTdK+aYoJH+UPOuUEm5
NHt3SHUs4puNMvK1P7GC18cbkx/HuR7upxaFo5sawy/sWwtm6X/WR3BCt+GVHHM4
+d1BLnF+QKonzoWJmx0aFAIVhKzuKwLapWvZeO9Bl9rn72YHTuZv63QW+uSyIgUv
3OYURRHGp1NUoDojJYtXuMkCYdFF1v3eUmO6sr0EPOmvEkBMR7mkzr2fjZm7JMkY
sI0IorvTA7NSR1V3mSrLDL47j04mTFA9tsoIC0m6WuJqDISIm4nYSdPSi3jRVwt/
AFn1xsuhRoyh3OR3M1GFlgLARwESfY7hF804fF88rWk/T1KQKTnmoArRt8xqUejv
Xm8TRXXoYABA8hi3A56jCil113chs89A/RSsAWEAmp5AskCGry3a/eH4qAx+RX8U
bb4NQEMY1sJgKa+5Pxi0RA4U3DHEvRswn6o0BYizJwTNspLYI0p1jFomdZ2r7Ddj
eGAvLPbOhaSAOEtxRvUfD8tcTlLErIia+Cr4NZbMfK6Bs/XJ5EiJvqo2iuen2017
9kRMolSj0s/U4XnCF7iC1AJF/QwZsVJJDwIVvHirRLc3o7qvU3NI2uo7yBzduHoE
ZFUgUEhcZz3aDLZPQFOocor5vm0SmSH+n3Dl5YbTjiXRkV/jXn4HfZRUlKqpSAck
iMMndcmYuZWQEXJeHBdpGwG8G6U7FH9ELnmoA0+all4tO/wVeLMR9tT9gtz2Fmya
bcB8jCKEvJManD75vcvbm7F0H2U/RSpoAbzFciAeasvYPhk3Vno38QbPOmNdpc7P
reWzx2gE2Qx4y6CRwTTrqQnXcQXaD6fw41Vzp/XK6QqtrUn+afnePPtaUqMhr6Pl
7tVwxDRiDUNGxgGmulW/UCBNtX7aeNF/NuLIsva1KsaTXLu7PglXj8b0VO72ykv5
brS0DRSxdr/qzFUeAfI7Xtw3tJsztNWYDQQHKHl/bD53yX/Sxn9C1PMQixKfAw5d
UBndyxp4tRVwS23bKVg9iCD06Nh2f8HkRDKyWtDgfsYk7CS5U8u3WUM5UUIqq3P3
2+jgsX2kU6s76wpIcgZZCNpPsjWFzjZg71jq+r5jObTkIx1llZCpPlycQADqv0YZ
ZkBP3eFdhGvMUKv2bbi50FLVcdxEA4k6Dm4v296sJyhnrdhmM8MTKU6JrHx+G+tV
vGyU+pTEgAaF3lhH+VT6tgsZmFL6hcezmIvPLDVT9pWxBfC+GLRg3z8jM3NaF6rg
9peWMBTIdMIDZXltarxUh4lf0Xmtqnxfd4J8OTERSb0s7kBMGAgR2HzBS89NKgRc
iwQbMtgmU2FGjhhs7wZGK8/RRqQ3GDdo0LlcmHUyvOfiMOTewFxvSdGsbChdODW/
sSD4JzOcXw4esnHhGHN+H19mYk4Y3htv08XyQJozaUzJrZS3KZynsOYQGFjNJysi
u9PdMoRB86GNCe4QFXeU3LJ+Ncii20DYbk2S10jR/fTiA6T5M6xnDohdWiP0DfVJ
nqd/QFDJPXylO8BlehB6fd1+OT0LR3uEFBU9kAWPKquMC5bBvlO0yC/ifvVkQ1TE
BbiejVi+Bh1i6NNzgWiZ2FWhPGolw+dJV+VYP5QLHKA+x+NlLew1fprlpir9DuR3
dJFvgpoddklGwLvigfEPHDl7+j93y+MoOBkvevXrz1dhFtMwOOL90gE475pFdEH1
LNkbcTK4okZcBAV0hoEaDa7uS2/mhjfUIoy2jC08Tp1bRrPz33Atjflb/fu/A4yF
1jaXmbN/kjFnB4p2WKq1zr8Wp8bC6gnvFuHibhZOvWZM7brsMBXP7xJJXKVbROpT
oohuBJB2sHM4svc/kblXeXKGjftPtq+fMth/Xj2mfGbY3agI9FOuT5ZMiXPyOf9Z
64HJzsO+dcopyj3pEgh8VP0MbuYxBFWWeWZ/qgSr+pOfbixjXxwOmg+CocM5bB+Q
cszwQ267Z0WLMMzeqsP+g50K3eTAnW9i/4jOvvsCuBcA0FQbCbl3MxVfTl+iU44V
spHQePzDpzmow+LUcQ9f89Ty6S1SF1R7dwqJfIgFDf64Sfs/CV10SlJ74oC90H3X
RJygKr9KwZj98W+9f8F6ZkKzHPdaYQz5vM1Hh5UhISQjMzfmn62daV9SSsGdwJq7
lG7wxDFbJ6AXZmWsVnlFhWCBqRRAGbuJfw0hnoL+7PKcmjL3nWRNNLjMSluaPt6u
M0d1hfUB4IgoFbT3qMVadS2bXXUdYZjFFcaGKbZyPrf9nS0Rh7wuzO1KdGqBXZz8
+zeMPYuyV2dsWoxkzdDfYxWvBqLLZR0irT1Yi/IZF1Ep12HmI3kwM/Sq8p8XJWPg
VL3dW7rnREf5TC6niLjYC6AdO1ZRfH3rMw4hRXoXVyOcDVgMzMC7b7CDXrlDrhFH
65ZOeGNu/SSVLDdV/+e3uTqfsGyzxwWoFZX5tTMkKGQEdw6ml5byLWbJo5kATgxG
cap1Jz6QVzaNv3wT5cMVthRnVOtSabbykbYp+o2dW9f/DSC5TZQHpbCT5FznzCOH
2kGgu4ifAD1mXh9rLH9Bxvrg27Ku3kWH3YIs3qsn9jzr0S8dx1tCDpLgay936aCJ
CTR5T+bKWPaUcc37CXprlUN1D6tE7w8mtXTNSDYSh0fXzWMSmCbmyyglHB24DvI2
LTQAsWZvBexoHz5qRUmZXgjAe2yBloAAZcUPKCaV7ik471Rxx2NVSE7Bdh6ejuYD
DCze98kpSIGxSHTX14jTn8fa0MglCyYVuJvmBdE/WixjQgPNxPzBgZBw2aeOXuQF
A9dIRdVAlNFLC5XDpos7qS5kBRmYtmttEI+FTL3iLD+5bwuOtqd9wBhZUwJmRFW2
YN3QJ/x4HlgZIWzzCpIP/ZraH+eaaZU0XhaQZYJXNSYzox41fCPHTEjh3eWVACBD
BKbpm/BmfuKhojO87QxyyscPXG9Noe37pkRboPnJrPZ/RdqxNlmK0pTnKZ1td3rm
+dgg3eEqkPqLb6qZTLqQMrkudOvBNFJHV01VDEiyB0chya0pwwpdOoCVzRXJrtuZ
tvccE7XRJJg7w45dvMC7iXASDCdvvXcJXdZeO9bhkSHzaVzmfXplkCC5FBZo+vmC
VWBevSKN75dz6w8JlMyFc/lWgS1ZtVsjDqmtAlgvbuZNQxFclW2iEHFtjIJJhEB/
kKfAyK2H2SSsmzAbL+4oH04fJMY/4WycP9eRfZXK6YSWDXoxjSzO+yya423OJ4wB
5O1Y6AYBK3sDn0+xBrMTFvifVyMFr2w6e+12lg8TAFgQClv4kQ8LIqvfw8/ZTrtk
JE27Y+PiRjLc0pKPmYbaoWwM80BTBPToG8XS6pzQw3GaK+651vczVNdzKQqwkUg3
zuED/ng+hpunIcwCEoF3t2b7A8YCynA6KIsxTW1j6H8yQy0dEQFBXWrit6ttWtjK
G2CV9cx+nTonG3KZtUh0zcz6gJ4/tRrBofz7cxKnt+w8dQ4n3PLsU4wDn18bJ8i2
5Jw8WZL60a3Ln49xQpvWp3DW504eUQ4NapdfPcgm5eOnBAk3xchIgx2iusrtw59B
1cku/N4KZc58kn6It50HLOsoriEjAMvvprZCIA6Z/pnRyG5MbNil9qfAxculnwhK
w6VB8qLuhMOJg7tEOWioqemqBT3IRYq3BcdrL/fThRREkE5AtahSpbGvFe0L2QKM
QLY9FgluTmX5l8RACu0UveC4SnHYFasO/t2AlA3KC8I19QCDWRyjIc2dVYkf0agI
VHel0dYHzky4xAWM+fNLYL1FH0PdRtyGi2/kBj00sWMqhYlYJv8KEkq0/hMf72Ai
FT7kM4IU/EDq735NT/47Ws3qWZT8P2lY6G8fKktgjPc4qoCBMI9Rj1LNH4/DUAg2
oOzI4dyFnRCYdJUDD/HfcIku9l1jwV09QuwTA6NZ90ysca1xM/M6Nw74r15lW0eu
ivFJuCkCaQVTgvxjCgEZgLBHQ0Vm5eLiHVxOubAeQdyhjLsixxje4938Xk4VAIPL
+81qjvDJwpU9kKSU4fOpRuRw8rNEzvzOhdi6r/JybKu/6eAWpzvt4eZl8eSOI4sE
Qmh4E0cCUiNc9zwaXlQT3irhp8oJ0TbCttcdr38VuMmwreDUb35vRsxTjxFk7rCH
tXrTrAVrnFq6HPh903biPvN+BBxmAkp1DeyzsBn3yfQ5YTTIwpIG1iXnA0XPOFWv
lhwRMQJfmAAUxaPFajCXAPcg0r9IU3W5amt5VPB+Zp2QIMhL2abUesEHBnl5K77N
5NrQWKmJAyfxj8e0ESQid/GpbZ71SCk3kYEPOCV+DFJ9vbyKEvLCB6l7W+hezxW3
HIsXi13EeDJLH0siSVnsNdC1KdOK5zoM9GcQM3+YElBO/1zsO/rFuKfcgPmF4yf0
5AoLlXc86c9a57qx7hJB1lTv6xpTh1wsfrTwk9RhiQhU9Iq5wD9duamjGzZ92nu7
MOCRDbPb97erIpfA+ZGQ9yz9qZi1Ke95S8xpVRacbAyLIC9+EeUUDGKf8lUiQh+D
invRutCAKS087vKcMbhK7iyXRsvDwKzdz9Im6+2OD9O1Q8mEZEvaERBJeeINAols
bNLuL4jo3qsO3mtm4o1faEGAJq2mOvl69nfdLDYdET52m60tgFYIXTG//JXw6djr
2VQzqrigesZEIW3iCQsxkzS5wwR+p8iURSmNXWdbcafqYke43+XF54llFs3LOk4G
QhSm2o/Ye/O6yYdSdoGmhjxKappyUv0D5iQ9q7ErRc0OFyVlxxbfx37IxRtCrp6O
8MIyn7SqWa3vtZyFSCCuTXtIg16u2A93CX2C2iUk6U4ZsZxLBYFwwiPM9Ecgqeuo
ICDUN1lzO08HsBprNuF9lve1VQC9qgpTJqdDcrL3y0bPmWl5mXH+s4G2283+sRxg
/R4sotUTZ3RiPMTSjNesB0mXYEJxbgFYCpmMpuEn0ChT66Nk4ZCOdZePiZY2wvdF
3ZMCtcWAv9mxo91MloPHesxUZhl07pT/17JsockBlSp+KVLQoJI3gvIPFmj2zsDd
1kl4QE1XD6yX86DunPuGdr8dHp19sA4Iar1G7/PkZ+Hj4NBKl6D3jhJvejV4YQtP
KRj04mXrQX5GRGGrKz+k4+S5/FHNPcAWw0aA5BZD33YacX+NQFa9EbQSI6TnlJVH
mVe7cmR5LMyHY211D0Js+3+aAxirLyDPug5MgaCvZhahrz/PrOrjLsrHnHVyA2Ut
qpMGfb9Y6vlaljf80YQX14Nr6Mp6aNva8P22cR8izHfWMAM1S3feSlBXttKnzDAq
fCQXcO1x+YfmZfsQ8POEZey8PjHKqppxbz1zUPylwUy8sikJfupEhlIOHybAt2qn
y1kO7xUAjwnKMaJNtKumQzR9GJs1cmeIr6PtJ8j1ZucuLKykneQg3vkB/qGedbtw
BB4fIwCdn84fhqcSWiyi0fQvdumnUCNEJxK+iQPygE9eL94cQC8Q743KgWwsEh3k
kMwju8aFyd3wykBKNvcMaEVYZ0srWwNL6c7drHsFdIULwrUL3pvLU8KrB/cO1njS
W4/c4oVj430jYpWpeIvw3rrl95NxXqOs+oYQIHtHwWAu72rLqzYPLqb4WMB6lF+M
EvS3qzw1POAFfKEPVZpn7lZK4jH1ubwG3cgJgViKdn/qOBH5r3fqBNfoIi8slvPR
BrHO/+ivh2JGRDjyfOIwzuAz0Gdyy49rKXlxFDxNJjh+AB3j39d6fYe8gXBD8jyx
ABjrSJS14NOW3xaUYTOVob1G6rdn5OwvmmqZtXlqsnWLiayrTXOVHSmEHcwsJDKW
fvci3tqgUs+/gS7uoiwUR1Q+22ymbOVm7I4alIIqpp+zBPLfWT2m5IcR2B0D0InH
I8km8+tfy1Vg0fT3xqFPTadW2bkW1LJBUbAMjCrfY4D7c/lb+dThxPRfmWtI4NvG
YWzguvT0bFWPQz0rgKWj7pRmk6uh2BnTyP3e58TqJo3wU5AHZR1iFixc2tH26gM4
c400dOt3fpdSEu2PgBbZ9N0z9pp89iOgQYQElIBSbDjcMJc6qLK6c+QzR9Wtp8sM
NYVnUcBe3OZBoENMitpi/my5mns/O7UK++7gnV7viEF7kM0i4S5EwcFsZdayh2Yl
eGFzBt3tOWZVuCNir+IYUKKmfUnGGKv/T8ymQ3t/bSZl/jYJqqPLlRXa7vEvpVxY
6d7uOeKlfi4szl/VkdNrQMppBTh+1RSbsrMU7ecpHtLqLi/j0FMX5ScgfLmK1GHH
gVYl49M1Vzh/UskVaaN+SPtcNj6sFr4F4ecTbgpV/JxAM52rFPzV/rkeWLIKkU2u
d5B3cuctORmx2DJgk0dJqv3hFzKESXTNdKLliFT1Y5nfYaDMryfaCg4TAJbQXEBY
6W3vYyg1vYyouM1nk/Hnh3ZARfD1tsMdtvAJ5ohGAaBBYIWIPnqhfsyxosljlb28
OYQ1hIm8v3mKDteI2QuLusYmjbIb/Sg41JgDiCRoMvsOu44gmccm5b6uETGFCyAR
PnTKyl6EKXyw5hxbVOIrOohORHiozwUGy3XzPb/AZz8mtuuNKRC/BFw6NdRIfmdq
BWm4qNf6xPvnn9mqxvXQhyziau2jlgFIpPCGLsHEZkJWsXz3rUXuWg/ZyZkvxd9H
AruM9iRr4wiGKZBzqbeiTi1PRtJBLqkAsD9WgLVbLWoFU4kOQpZGjw6xJxrjFC1v
Et1+NnhFiRvxnrnF5DolfWqxCX7eOoF6B7oYiM0d6fvnGXbfF/6JZ0z37mEGStGs
alLx287oy5+K9Om0FIS16aANmJLrxruxnRtmjtC950f16lpuzqffsMpkxDfQCbYx
fahq8RRLWiCAlW9rXd31Fq/uuk1LtXmu0E4QKnjmiO3xR1qEzp6PjGd8ls2j5FiP
ct8+8boewhU/sWZamGteoQ6leSh4ETPEqhj9q3F5PXv+Mkfz2T8IzD07dvoLumiZ
MMvyHF2g0e5ttKRNFlX5LPQLZtidLW9uTWkHdlG+HGSYxCGvrMdTNkxhb+YAuS6g
liV5OiPlzwCwscmpYUEMjWY36MZJr4T4FxCxZIMIV+E5TxrH2ekkn/q2FbvDKp9x
yb/2s9wFm17LO3a/J9NtOPdI5U6q0oKvP8QLZRREJHNuVrcwLTlqqFBrRtidxiXm
vSv9pUKE0LMNSssJVOinJgTNCrfMgjwgbi3zLavaoSIFS/SpDNWRvOaNppdRQsFg
rZ6wIlrJ5qlkrWP2zXcvXIaEEAgbxz36esMgTQCEA1KuiTvhra795u1vSRrOY/qy
ZI71tu8r4/Mczf2r/0WAesEvBfIe5G6N18qmVtUHnMzRgY3ln2NoQvsMrHbYu1Rh
KJYqNzQRLk91AVNPczhjDonPao6y6XFWWT06ZEAtBrak2qQtjBoVrFjbQj4B8GMz
iSekcJI8m0wcFpDEvpAZQqYOyBh8Gf20DndXvvFWThYxKyY62CsrQlhiSjpDNiK8
20xgC64x8HBk0I5CKnh9Exb2/Myu1fCDlnDfhoHMSYDmXxjhS9vMyhUcH/JqpWGb
R7U5MRjAAdyQmaSRB9cFp5Wdt9DwCDukPy3iS6rM6FYw6nDnCr50nsjEAGyjedgb
Uowo7mP430HXDbzgri5VW6imw1NC2CrPvagtt6ALAnVjIET8ke10UaWU4BfcODXu
ezXpyv1dead2baQi3r8eUSvvB6atx9D5LcZjPG6n+7gk8iHW65mlHtGOpfEUNuRU
2Pey9pGqjzSz6JNYI2mUgTkWlPtjfpH0KJUxnikWHi4D0uMY/gnKcp8uGoDtOatU
cDPBvJKDgc/NwgCAF00P0OJDMCqpbazi4EikKM2YHgOH6BFBbaYUpmRd8/y6dL3l
iiGR7s7C/FxikHewE6LmJfHrUCH9u5s1NwY86x2X1STP1qAH4VFfmXAamavV7kL6
33jsJvIN6yw+nWyyiQj3Q4fjxODxM4pJGlJ7XYOHRLOSLPbIuyV3xPLIKSSeTADy
hqIykrx1etb1KAAE5IZzhsv+u/Rf6TJuMy0Y4isLIwFq3F4EFoHcdjnxMlftXre0
z8rbjPoDrms5kVtD8aFhcKrUhWWEtxozSgt+lEbSJsZKPlIKYWpYCFfKn8KaGIui
XaEwHxxofTSmGiDzJidP2TXPnl4kDLAYV3bvBc1ZgC7xKLc9hFKAzpCOaOrZqDmP
VXmS6CoYaHt+q0YeFAW0q7vkUkuuN9s949J3PkVkRXSQ1xI+KIr7ZnQMrSQ5k0tz
gJEg3FjUM0Kd3KnQoVL0ZVfCtowHrLu4luiGGaC2Rzw9DBfRk5Vi69ToZjIiMx/r
RHBmgVEV9d8WJXKicdbfnM2YehSQaB3OZLR6TkK/3p6LkjWZcdYwWrszBsN4SbTl
WgS0QoGN/49QND2uWQM4iNOzN+bAmTef9HR201mcsi/ifpDawl+XS3JEcEHDa2pw
NSZcJ7APK2x0/JOPhvxOEE+6mbjYr+BBjqZqnZuw+PlrCG0iQxypEiljN3YuPPrP
fZ+VsxOBafUyVKHpPn9ONeFtxQ+fZ0g02JagQwceU/gvWVhzFeloEFZ/xJtSXKPK
JWtUrigEIyh+wzLh+pZbhMMxkJbVBXSi7VwkjKb80K/h8Jbdrg7OzSLk1IzmYZDY
qHhgciktdOVGJAYvZEri27tX5EsC+9jGBdRQt66EqrdMrMixIN0vFVb6PDE7IFls
ys8nBr2dE0cyU2Stml11ZWKZ5uVAyubPenafI3htmF4gpJCVg3fJh7E+DVRIGKZM
i2gK8nPKBE6+//Tz03ssHOYMin+6JmeIvR+IbB5+M5mFJ/lrGuCFhKB79poC3lHL
+5Ch3dQyuo+S1qKsEkVh9IQ9hGTXAaYIp3+lvhStsaaR9p7D1qoy4SWrZjzZ8qJw
azN1H+L4vpABVqVhh6iqHIw3KYiDvZORsMbZvI9yELDY/+xGlxrBu2yUfjaIu4m9
WYHVBTF3BF7coKWJwM/DwWEYcVViCHG0MZcQrWkpgNaHYcSqZq3Sdihj5fq+05nZ
sK5TmvfH+BRNMV1imLINxa+i20qMkXuN8IClLwopH3DGy1MH64EqMwcrShJoU9fL
KL25zn/W2BB1w2AYg8lOqwYSWto3nyMr5j0lgypKP2S2KnwzFNY9rhGEzkk92R7X
vF1z8rQNabukW3EmdE4bidqhXJz21pEtwyXAa8QLegl7EarNG7gkqec7ZSsKrVr5
f8DZek0n3sAotmqn1UqUg3nC8tH7MMaZdFL9P+6TEjNiDBZIgjjy8zTMsyioMbLk
sMkZsynQi1Ea8cVWBQ2bMZKH5NlDMV91Fn1yl9+zOVUlLFEQjTViUcP0glzmlcb3
EzsLCyicjWvjze7UMjpffwCSTqenkQceGBExzld22SqBfIddB1F5SfF9DxhBc8Ac
ZDFHUBw+kif6c5vFM34Uyi9FOro2k9Dk7gD4dU3GAZfF59owVCkOekAfcZsh2JLy
eG40K6/uun3RWU0VhpRJsXzxUEobzAGz1+uv5UBavALo6XxGCYsQZpQfBHiUMl8h
uYmRIxZWlP1WLfF7yvDQC6vgq2GEbjNb3IO05/wS4/3CJqOoNKw1pQnjUXmXgEYR
OIk9ho0RdJ19bRY3r2Z3SD5prIUai1BFvwmzLEynfn2JPbsraOgLczyP0dgXaNDk
/w3FMpZwUawc7tyzZQJYAow74zgg2sg6T6MwCQVmwISh13prEO/ikshtDnw70ABB
T1NGPppoMUUYv9hHzYd8Po5CAB9cxiijAZuHipdf3uX4Rojx5MQ0tbpKq8B8bc4F
CEZRSgRZ5YTXSfhEUxfT0lNZloXRdgjWW9A/bWxMmOFG9+5WsciKWfDOGZcQt+6h
eHzDtPAQANa06vAQDZWb2cE6yuvCKYtqwyrRY/F5lJg+1Uolvu1INiIAg3yoaWnC
Z20A6CERbhVor0vmh7mOKFnTmrZSoZqrd6KF/dGkQtGNyGDy+2/gq7Ds2axY4gmU
1wqVUGzqNR4h56cwEN93BrRfCj1LPmQ/01da/JFjy4QT2BcItPuER9W4oGFsqGXl
5bbYd5AGxqRdMdCNacbMZdHK4dnWOobE0TPghcR5V3n56jiWgz2Pxt2iRdPRzinF
hS1ZKpJgYgqxuED99+g3eoeq6OW44nG9UWlwEHMC3h/xhH/nt9hnFZNty22kKTLD
QbxTEN/zMHiG/mCeaWo203No2QnLFxhoHVknDURPxIk95WFDKoedF4JDxjZzvJAo
TQ62O/NcCsacJwrQSMEkq+0ggLERSkCs4nnrpNyrEC/i22hAAVbkJB4Sl5fQaQJ5
8Gr2GFttU3u3IyABRWxESRI3VwoaP4et9fG9umSODn5X8kV4uZB9eRHutzod9QZK
W0Mz++1zBL4iXjWzaEkSztq6dbEa6wnenotfutUUF4Dkczc9Pr8DomUqjZkxSu/L
LBipsCM3i+TSvVQs+A4VoFcRmszkf2ZR8dGOvGpQiaGxP92H4zuH0YG2mBHYN09D
J/olNOZgghd+iWPkDNtKeqO7fI2xdjhyN3ahlizb+UHZ1tqjuT8j9tsJSnMue7dT
TVbzWh2OUu3R9NbOU5MIJXhA1HoFYKWRmv3LLz1v0/6iDsgIqueFv//vKsGWXPod
X0yBjEI99z0ladYcI23lCBFbdhwCkS2NrWMzPQ4JyM/FFHaVV/pAYk/WAfpp55ms
xvCJYEy1ikOTSObYlAtMf9TpDyxnS7mvI881rJfHdIebcW0XlNnl5ful+gWi27ce
IHgq9hTjivf6OFOtJEe7Zr7JVm6W+od0H4dvsrU/H7RUZW7okv1TaGcmcVQzjl++
7aEClWgpg0xC6ao9Ayyt23TPqYtEraN034iMG2Y65ICQ8pNE0kfhzM5iOJyQnIz7
5OsYZOSkIfg726pDK193lMLjZ9Q/09f0lLil2OQg3xVNvzAKTb8dFYgUQWkTVTMY
s1aH1L1p1tzU9Soz6dzAIzybFftLZuUwrt5mEfVfSYM1Kpx0kJgTFFCim0NP6U1+
U11FQyFQbZfeT6hecOvv24UP1DzVucZqPX0qBqbm1t2tlRZtbzHVI9LBFVH41tPR
sYWcFKqClMhaKvENmX6Bf2eXJZq/0w73l/uGF7ohcaCNHQn4sg1wcfsLWrnN3Y1r
5f3WoXbzh+Aou5eBBvETLkeCmt/sKtk3v0DrmvyjklAqCAxR1AoXGmBKEbkfLNEl
MoS+cdgnZPEJRyvTJLEdDTbOUPzCsnA4IIVRYHKyTceKzKrdc7vDCHe8ZBCYtTsp
akks4QFuS9vuJZZub8ekNFAFa5qUvOTSPNuAbso7Gr52BaEZOGmN3cZzO0bj0cto
pATrPyOZUSl025Bqm2Slrn9uIyrhuuMDAY/HY01QPKPwjMHuT4IH4zDV3ZJfDLcl
P0biO2bcVmv6cUCYwLq5DYMeq+qA2Yq5xoP9tpC8SvMuqmm0sOBvdXpKnTnT8Drj
IquQMOEifpfV9LbJJmOqr+wSCoO/7qBpWoeyqErMrkzEz/VjULFpwlOjIIB57QBO
S/CMl5l7tlSeF5uYfkWI6SQTK/thYqtgIsujrMdneN/4BGjhsFIp9B5AL/r1CCPu
zuu3Ol4RCXq0bc++ghZEwCtIDi8ZAP5ixtDbbU/5NJPauo5B84wrF319aws8PoTC
Zlv4fclt0j+pT6rVjLGvUzAaodjG/+q/6zNWGLwHjB8ivAot1NiO+xMRxb7eldaQ
BC40WMXPN/WsLi3jltAQzy1lHSb1Lh0nsTbAQNysR+CmVLxvvBmfkFFNvRgcmNXk
5wSN+yHweS7YqGsGTWoE8qC1No1yxQaJTSOYX5YG7NFWCkjjoWu8egSkMUBhIHOO
9KRv795bnJ6UFzLryZHVEQkYjngeWzRCaicnLtYhC5O9PLCHg/KVEq5zNAnEA0hf
21pe4bPDEQlirFbFxVWiJT/u0fljT78HbS/peny7wLsA9P+5zkc9O9M4ooU7h2Ax
qgA/UIfJra0e2qlsiiHTn9vQG76UI5HGkgQBSY6EAbyYOENmSuJt/lMaX91H/+mw
sy8c96NIIbJO7QoFu1t/+NFAQPnNoeM0aC7sfZXcBS8xdHvEHtuWKleg/BA2pFVf
d1XhaJBEtsaa14IPuYW8EsYLHJ/LI69L0A5Ng4eXnJBC8IlG8xm1Wl+dwOZk/koc
x6bgVYdDvC3vkdmMBI6ifYkaUY7j1KF6VQ2/TdD4JNo0jY3SHDRgFeOEzIy4P67c
LgFI3UGHaqQS09su/KwHyjhLDwh7BgdvlFDlkMB6vowKzEMgCXgfT7B5ZNH2NqgZ
hxgoXxdlpa7Vz3DoIkh9fkpTfgFih4xMNEfemhvUZiklKURdoh21wYXwJaI4k3Or
U6r9me1/O7IC0SCbpaOGnZXPajSe5vvW7kFze0dJGouN3KEGM6Pm/Nd/Wpa/HFYo
WTzkcMxnNeBPeCgOF40SBAGXgaygvKdO306JGsqp0+9zMlXIzlC9SqBQoGuiILW7
MLfim/KAhsJ7VmfvMXTI8bF2vxGZ21zCKST5sWA9duOKlWIKjaHqxyXj6NQhkIR3
HTPAOX92dZ7ldBbPdjBfuE2Nyespr1m11CdMg2vh2ENrGQhYruddChGgGN9u420D
icgBPrOhPvamkLfZFNd4VALiPL9YRwkONOg9GmnmviyULmwm0OIXmow97v+zMnZi
ikZBd7Irct4rjuRtoIZSpoxjtSuzCyZPx5NKMxEvZmqhhdMKFaDrtch2Z4fiAaKO
aQxpz/bBd/iUFPnEns1Li+P1YIaJ/khbuDd4kS1myruVc6Xw2AnDp9vDZ+THHq2g
/czHCddRh6u/kChX9vUb6czpL9Uji7f+mDqPRvJjA14tkUcJN8yHEMKaWIjmYBHf
XpWjIT0jiKf/GJeXYPdI/vGWxYVBAMoL0/kLuc7gpFj46wlbDxEyGoan+8v9V12m
gRPZ5O+4FN3xQZXAbyjhOwJGZ7Ng1nXvDAWYaijFHklYJoS+Tx3LJeM8We7juJh3
HL73xenYOTu/EiZ2bCThUATM36upeHchf74Z1sUHSJUKNoJUoaOQvjKh7wQQCf2A
sY/GZRXq60qT3XAH1NvAt/jgwojB5787e6QV3ghCnfQt7i4IfmnBaWXrIq5kdAVO
GLdr6Smo3+6LEaCFgsEkcwil4yMw/sYTXKJb4MPJqX5FD8QvhxaI4pMTMUg2pBj6
P+yxwh982sWHOa6iVBk+UFVigN8hX0VDl8f6VMyskQeaBnyhw4GNklNRMioLb+DO
b/xKix2uix7/2eJnVTSW2fKh6IEOg26GL++mQoiuvyjWy8HaBu+H5gHBjhZWRWd/
lqj2kCMTzaoO8h9VIa+KyS6cVrEn+zC6Bl/MmPV49Jzb+04DFpC+GysuuN9Lr5Za
3Sg+xiL+9TAMPIW+fshMKKYOlHhI498DRmtfMMFVW3UiV+EhC9TPg2zf/R+bh6sL
oZwQTTIMdNk8vmDjdSTFtSUkXZyMCJkxB59JmqatYYq44FJlwjasf9be4I9ZthpN
dN6qXlmkzvnQTX3Wkz/2ROHcSaJivVDlV+99LyjaGnTIY4rtuCxNfUU2+G6M4Cx/
Un5cC6BtGON7OgecNCc2QMCOFoPVefnmtHXMTvhDrot0eEufE+D/cFr7FxJ31aOt
odRav0CoCHfLHUZQynqmgJWOeDNjG988/QmiIzYwttLj9nARYfKy3EEvOtS/7dXE
yZr4stW8Phg86X8aN4SmQLHFcgCokOQHEbHbSZIgEfxajCmQDkK/ps3nJl1iNFvB
OK27x/LmBoFi+nBEvLUsjhm/sVDAAPRClEF/R1+aoXR1BtsF/N1EViaI9Ngey4wp
/GyM1L9FYx7o8GUPZrMqmpH+fv7yeeBhe2QI8Nbv3dyezXuSTJr7/im4Dn1wYKV4
BUu4yLjaek2rAcNWMyjHaojeAJ2o3raFBGrE6+kolIAJfe+9tWJEbF76zQuWreGS
Tydtfz6pzkLZei/90Ci43yoWtSvelKQylbw0fzU1JRnYxDN44qmdXb4DatNN1rN+
/vLloY3qMdGcvsFxXwqstj/2mlhkK+eDjEiXhJA6SuJgfSGR7V1OH29vMtFE1tvs
KE9FMLL281q64IplrrilFVuG2rV/oTQ4B4xecs6K6zN1pniHdXsYVvUoRoCglaN9
VenL4nEtd5UrAPkMnZwbO8uzuxmNUTCQsB3CiW32nZ0X8AjK/zhGY9s27WjIu2nC
5maU2NeggQNCdesqWjHHcII+EP7CvbivxGV4yXNyJQfqCiNa17DbCMRS3VzrUjq0
tJu9Ys/s3BiKSVmytfULM1VwxRW5YlsRejzLoouKrrLV8+Rt/ekVww6s7lYEU9MR
rd9oADyIvl8vRi29OLNtOZjtv6woCRYHXJW/PNT+7d9b4E6qb/ZVNb3HXnWsnv5M
+zd0veOgoAADaTJRvpz2mk+SNWGTJCL0z78UzzhTwtHW9vtN7kE162/B68Vvb514
EEMOclSui8ciHAYT7qToiLsGnzU7mNp6kmU8hn0M0lUgvGPzPziyPQryTHiPhujI
jpe1oLObzIBhvfzQK7PLu9Eqg7ZJ9/YYpTN7MaWS0oS+ewo06G0d7qcy/ZTHiTIG
8tqoW9c5mr00HV/TVloZ1gYQFxHmOqlIrH6QJHM/E7/WULncE4OlUOnEDJwJQDm8
BQYdOYU/K1Md14F+M0nYDDJsFtsErQvfJQ/gKsGgWyh473Rt8GWRjxNoZHcy57OO
ObnvXAGUWCe7wGyOrlXqCy8OZuCvmXycyR60JFUf7hPfOHtzwC0b1NRkst5QhVGO
UFpuI0UXIgU6M4ON1BPbuxmvHzlIi17fAa1wuGG6Xuf2Qe0T6nfIXcQD3tihwWzz
Z1/c49VWjwQYo60+toEjwJmOLtJu9hqv97P3WtPtgB26hafmRe92tUGsz2mCDA3W
QSMcLysZbtx77+aCWJTaFvx4EDxJYuFVAkbajhHdbzhGE80vqB1TN5nC6ZdKEWrS
wAbavVX5+newjTjnHdBTOflon+LYQs9/eDvt3skVyR4YjPUUX6BCnf0QANyJg/4I
/DAl2NTU7VBLG67XAr9ci/H+V78GR/TNvZzfVL8a4CqQsfuxEt12GBPCSOfYu9OG
P311zXdRwTivJxOvfr2MYdlrZ4bDlwaiiGzNwff2ziYwuP671rzkrk7LzkV+r/s8
1WrMOGkTSq5Ig9RMsY9aTOwFxoanVTomhXacIHcBbNXIcGNavbpTDHrSgd6P+egV
zga/v+j5cHWi1y9iSl01yicZnOdcAv3pZ/nWTaYmMnKcXh/6MGaewJqQmeOuxgay
yFEpuCYy4FCbtLO+gCNFKK5nfmRVW87s/xLMNS0L2v+uoNS5r7wWQfKtoDX5Nt9X
f91uwFjE7lgqtnBHCmA5DSygkd1daslSQ7e1a6SldccNvKYSFaJ6AfWWLIAAiKln
Qm1m+0C9z9UwCWEVg+wwG098WpMt2OivnHUZuQj71d3YnK/VKqYFXmVCsvjiNlAT
JQMYZjNAJde7bObrzDYE4kOarkOAnjVtdjWUJxna7tnRhsntK/ltZ25zo+3mQfM9
s+Zf+cBBOOlrTpcjXAbmBbz5VFHLLoCUft1GlHFsYb/liqUGwNACIZ7iLpC5NNwS
Ehw8qw3hKM47JPuUefEro4DvLqsMSWzZPAx3qT2Rq2QW9Bm99AaUl/Eszu8OIwQA
6FY6CynWlYw0YRBBi2f2bOgmAByNuJEI4983Iw5KH1i3lyc+VjOBdEnsVdTQxC+m
fgDUkaK3QnA4D5ZZZYHJYOzOk3BbVG3ehewhQvweWXEi3TL1uj7wqvX1e6geKuT6
JjhOqSs17XVziwCbt8ox80XIRKUmIERlNewIZbhOkDOT0jxt4iOctE2CN+MXDhRS
LAZAtPKVOnaCn+EsGAGe3O5pvEitruxzNG4LIN6+c3jMnuhl6W+BdJQexSFU6s3V
S4LEOXszFG4NTdeXhNhpxwDG/R+uagFJvx4D4RfTOyhEX4F/kBklTW63yU44SK+s
Wg+fs3TvxDPcLi7QzwgA+B60RpoO5YZQz7hABuJCB4qObW26Ayj9/0jdAdHJA/9m
KjNQcYhf8kBibx8dws5u4IGJ4JMjwbXiFtiMXDoQIbC4rKcetT8EMDd3qYVWPtKZ
UYLI7hM+UHXUiQXG2bt4IOt0GMpmNbnHV7GNxAVHYEG/D1K/jY4KLGw6DT8hL7cv
56pug43TnReCChGzCCnQvIAmGLCVV8gqVST/ifl7f/oG1MZpeRM1hkiNJ+uYZXPc
5FgParkgmIdHSZX0mBSY+lHmysjCxssidJimO4tu5soQ482xBu03CCx+zMO65AyH
Ta9OzM7jePWu9XuIHjaYUWPLM8rghsiaaNE3S/2bmjsIHGdXt9HFSmuQ2Z85B+pH
1I7Z6O+1NKJwRcPHIpANIxU9YYuDARRNiKoAx7u6qwm4fQJ3XB3zKfeXYZfYMX+0
+JH6xJz5jcXkA3v3GAZhR4mHxdhMp8jEdU0IjlwL5iBCZxfj9/wc0+8BkBukmP81
m1qNNJFvDpeVe9KVvSTyHcLpD/goMvV7Z+t/rmyOt4qPIZFmYKrUGjLJY2vzkCTv
SthfCZBjLoyC/01Nk1rK9QuEkQTLE8PFUnHhrrzeWYsjvYGEFZuSPsAtgl3q8tgB
j6z6799JdAGXb7wQ4Qo1UbiXFIPRlJCuwMDe91KmMjBZ0Wlr3+iPrDsDZJGKtNVH
uKwwWWdPZKFtO+W1LlQmYlh2pHsfAfEvs/R8VBtvPTzyE5EGkOsEkT76sHSmJN8g
DtX6/Xo/qYtqreeer+g4ZvVDzsgDuRGYtKZcwllB8p1aX3tFVYhepmIXPIOc4xuC
4UtLK+f8PtOc1YHtz8OKJ2df2/Q6+0Wzm4/tRfHzQWnY30aeL5W89Z5DVUmLbD9E
OskRSiUgmkIMdfuK85NYktsiKaUNYvKmbubHry0iEN1VZLMHod0J3ReEa4y0Y0zc
rSGJVf9DkCCc9Ww8vm0V/bQ3EpPOUBitGH3+FjRI5PvygULReBS3YQt0nScuCtlf
ksscSREn6XPFwsVrmOkWIiGSkUxt6uEo/u6isUX+pR+B14+xoI01ZIY2Rj3Y0owY
lFLiyhoQbGqnOO9htfY+1veJYDj7SRFbAAdXgLUZQIBQ2F7IT5yehT2LmQ7thBHg
OOWUQkyyh1eCyjnsQ5mY+NjzW131ZtfBP+2h9M8HVueerJK9kgxy2wrKahonZ79k
htck/7THyH/Ul5LBIn35W2hvQhMt554N9z4mafkIR0GyCPWYEzVCBn9S+h+vDeGw
VBzFhP2amoNqYdkGquyc/IJeNdK+X0y8ujdYGBwcryoszNBGYz68zqw3VqFotoVu
79Rk+GtiP7Kfd8L6D4R5WozBX2JEIf18NeF8eZupu4kzHgX6wUifqNGtJ1hp17uC
RDKYd4u+88aGG/JI4fgLvfDhsFxezxna/Z0bSBlJR0IOnqc6MJtNXZH7PCAqGnZD
i5O4pB6N+fOHHCkWyVMeKPMj8pNwVIehOTtYlfiWT8jZRR896oxItvJ7YVPqGUQy
+ugbCOByR7/y9/xQ23P/aWEj6rPPz3UXbC/TVRCwTpWIw95os45TcDJgLsk8fXpV
AeV0zhCEOr8qkyAtuGXV3WkHch/HDeKRhe3MYHeMI2hXT3v5wVMLYl5gtzqGbF83
Yvf8+BexP6jaz783P9eKT7B050AKLn9CXR/BMCYhnFNJOif0JVDGYTo2VP4phS4c
+u4RX00sQZ596lWDg29vDWeKCRW9CReagtrmOFaNxgqoT8m2Uu0kYJk/aI5J7Pqp
1kr4S0oxcugXORdQzG/Q+fyi1ucGhlWzcfHo5jYIFoRVlTFrVMVtpZXeqgWQRDqs
0yLCQ7QOGzuj51BIknR8N6bgXR96oMGZoib9S6FRKOzBBVLNlW4WiK8ClVySji5A
FkNx6Ve3bhOlylcWSIU/iMHesyy6+RmHai/9YbuPP4GscSiqXyV2BZA2Rb1tMVSx
djxxOK5/uc+kFV5+Rw+nP3+NlIGwR2rb2LafyPvnP/FcCCEPlm1+1gqGp4VMEMAG
hHJPoKk9FuRncMFwnpyGeBIv8qbZj/u9MSy5pBLmqMUQ+N1+ShhqsQ/zaL0HNgWm
Cp2cVQLjf2NsSxwuT8fHvDM0gxnTQz9WOZorvotCAqVAKovgudIeJyvtkOIfILNW
jZrDiik+5lvB92yPEB7DddH1ebGL9G70Xo8PL7BAHQD419tYWLLsakFR5lDM9vJs
6OroIYosVBy+XRYAIGcazg2oRb7J3d7R5Fl0dUfqOlbPHaVlV+doEY6R9RSSExYu
z7ivVjy4tfprpzgR+gYlqZxN2KngWR2jsejN74XMP4EiLlmrURgvO1SjW/q6wHxi
PKa7EHctJyeEgR8LdaWoXNhiXRcoHulxasrb1BHRDLQI479WSk+S3Ey1OJFNLarF
BuQmUNH2jIHeQT467FXxDnTIyu+cWLdME5/OU1gdw26TIUUVaTpPyIbJmJf6dgUJ
K/01bAo1iRwtvnyTLe2hQ3fZfPCwXuhuMxAifvWdmeWKdL2ef68gwAhwss5mvulk
edsrcV5w1B8qEiXuoOkxq4NusoRBjxoYR7EaRMVA+h1TnvtTI2y4x5vlVX8JheTJ
Yj0fXW6tr32NOciTIU56+1P1FtZa/J0RmV6qhZrzFDg3bdcLm2tqxkd6CXxyOa2r
QkXxsxWu4YTHu0dC4GWLVINkA4uQVH1+lqkvXV5H5jSDvYud0+lWXDkqrHrdd7bz
yTfZWQeR1HbKaHk+DSrAtFl02fXva6cdqyz9v5ifflQQLDo+kC9uS2EYwD0WaLAL
oqS5vq8lQ3CQl6lbL6Ul02O/TElnyE3bILfCrCxEzqHLuuVG1/FVWEr7hiF0ds2n
hwVAoOYYKHRIP0DwgBI4sqk/Sm1rt8yH1JFKvv4gtrUQJCY7DpLNpQsJPluKBHka
0lvbdwAfClacVckFsBp2U/zPz1lllXXVUhyDqVXzxtTnqcr5mdvIOXcF/NUltgS6
ACNlX1o7XGXq5gn/Re7XH+HqAIdkyK43NOqdi1vpXdSTi6FLTL0EWqnje3J+kShm
TlU3qIlO4H675puREpDQdroRqAX+z4HpNZDGgLh63lnEJDFBdTvDGyXXBaNCFfG6
uoNMayCPmY2iit8oypne2xveLiT1r6etSWVrBsE3FGYjB6Z+K41I7dy0/uaLgJJc
zl9wrmqHd42p9pIr3JyZCj4syw/GVO78GG/DlNP/bsIGTEmn5w2/LqaNNdTqI7ZK
qTx6lY+AZhT3yuliyB7sNFSsCaO2oiez8eLYNa1m2BkBjeJQuf3iD1nA4yGCZ5ri
AyqyXRvv3x2NqGZgCsXdVR3osNpnUVOC/gjxTJekaI5WtKxUJIARVkLS18fqWrfs
dvAOB9ruV0meqkONK1kMCCNOp7Gi/50VQeSkUrruiafHuJTVHU6c72/F7ObjgPHP
1qAPWi0nkZva1uA65/KpXG3RJmGpuGp1npSgHQ3Iwmhnax2SflaL4uP2FXmgHfnL
bT83Uy78ZD8awTckGi2xf+agRqqxEE4OyFu3BXeDnJoejq978Hl7uuip7+PEkv4K
jkTDD3Rsxn7KAzt/417CjCeHHyz397983atdK2xScWYjLniGH+JYMRF26rLUvQuM
CMwLDgKxA2ypb5JNik/mM2GQPXkTKskiH72fWrDxtjsws3bnT7+hgFGEL19K4cR1
m9Oq50MVML79FMZd+PuQDqINXX1Q9vrfBR32EY+/dUezaXJlpJCEnbXpbLnjKDIw
ldgZXe/Nmoaeedi1+B2qVsVnm+SYscu69DTADWkowcLsOanDnZS3ok0szSYVSjFW
sE8YAWtqbjr0Nukieiu8iIjAgJZpaaQtH9NjGB8Q6kLXJwOvboROx86Ms7FptNm9
H24Y6X3nnM4SJOXT9TviAGJ4MXDXqhy8DKA7S19QaBpkbA0D8zbFOHcak6DcFZfY
7DiGr7ObEAFM34TDSzvwCfRjFXihfojkUEu8Uyy2lciAxHVHtY68oodNFvHN9Y3Q
0yLpkgpsZVIdU4Ypu5unled8W4sV3ErCY6I47QCBKlMGYoaj6jxdoxx1ADD/vSUT
T6gCjpKNP+3Xc7g9yvg2QZ3p2TiB35gFLL5Ote2vwnLI1zhy0iN+c+OdH7+Dtyhy
LggV+zMYwDbEASOc69PL4994jI3VZBNifr37c0pBNRKL1Bb+9N5YbdjgT8QBN4BS
kjoxD9c8l48KEa+QhuuOVKVsHnYfMRkuqipLKjVKqnfJTMfRQcWLrhaQYiCQxIFn
/sQx3VTlNXCLivQG9eZXD82WKwpylnYC83HC5pTrHqVDflKrXhgOSwA00D5gqtz7
est1mOXnv7mWperYHT1FkYSLWrBU1aVNErLJhM5ywqa2+4KgDWoVPdzQSAfbwqDK
zqgN+cLganWIup0kM9iibUbN0z/822W7KGgzClNvp4s3GOATDkxpWLHbVOUF5ulU
eMnxR3cKU4qzc9qPfmWBHjutPX/JNV4lIp8cWSAW8e8UhgKnjwnw6qNssB+iRxD2
fcRc8Sqj6mSqs/IIRJVeiXBPqUURZu1u45bfTSChfOdIlNea2CTe5VFvzhqJMqeB
NaGKhrGPK2B/kLGfnaBh4VolludjRVBOOXeQHLR3cPDRxb8g63STYfRszLhZRVNn
jAubROhiF2HuIW5+WYHqeEgNtlHnEKs2I+eDAIGEKb5NvaY6N7Hcuk7aWiXB9XpN
JAPFj18rh+QiS1Mp/jrxJ13EUlu6zj58IylCyDS2zIpKjO4CjOT7SU7OIW2h4TwJ
TzaBUqgQrTTX5n1H5zfbjZd3HqN/QCaFp8LxWPupIa2eZkJrOehUDwyFPaXg1eT7
HZatvQlgrjEpYwAbznD1v3F20qQ9viNY2+SXXD2csRn/ThSeaUNIqn+T++Z7JlAy
bzj/R83nwdQy9m7DATmkZRY0zNINlZfIKMUVs3mz0quheh6P2hTD0asKiXGTp0jg
l+pxqKdKywmG0mxkSJ5jbQ/xvR7JiUQ4eCVcn0I+R0S0pvdYCh6A8bmr14L4L/sP
KBWnzIN1aeHQMXlsn7FTCNEmcp/RYgG7TfzPM3A6NpIGv57oE3C5w2qmOEy3PQ2D
ShhkxD41xMEOatXcslvNEjBN5N01PPJMxbIun2uu/vS4ms2EQr5kUe1zv1jEwRLL
+f3ADZx0AmtX5OaEXJLBqOdMZTq/a9tMERX1RwlJa3FXtIbILy68IePuZqk9x8yd
s5dHYxeMyw3XFKeplq1e7THYCw5R42UXNcGMVmZqpCEZ21EO8+SbIhEPNZ3FjKoH
NTMu5a7XXZexEquXCUF6uzls9ejy28bvPlHR0UXPVPyGddDlR95z3ST9+mMluTgC
CCcKwnL3LNIiaXzSoUiXG19nVDKviQ0vZxwb1AVwx5n1eQTaNygNG6ju+npnFdKx
UuB5hFCLXQbiQtHmc6hl3YumBHg55Pu4gI7vPHAuoP9+mXAVmGqS5psFKemFdN54
6UfRqRVdyZh5KD2V1rTJy/xM+BNw8Dwa6YVxnSOC9QHyYM4nmy3AxCUEVaKl1Yr3
7+WWgYMnDYZo1G0mLLGIVSuBB4FPy2WHapGwLvhC1bOKr5dsoyVpMHDyyK0+Q/rS
qPGxd6S9/KojC6dBD+yOXEJWH85PGOIv3AmXa7XmjuirkpnfBQYoOQtBbaK1OBCQ
epVuuXf1I6Q0HU+jOq16QIKYEWgyPZJJP9yGwkjuYClE56FDp2AXFPHUQ8ddnjae
crjmIbAYhCtCzcMdSNdr08qtVF5NINSOmnxAvKIuytKiv8JSXCnupnOePquW5YdR
QA54n5vQBAY45CFsiPL6fmTOvR6L7jrSQ9ZNmd6uifC4qT54yIew2RX/57Hf7bIP
ytMrN+QsElFnFHMFJ+Q3F736ZHUQogvtXB6OCKXd00ahSDp8mhoOEjUd4leC7vAb
OJFeN2tzZXdkLOCzUWorhW9iFE3yE2/U3yG0tIctqwUHQ/P+XmG/8wDqku1VqEWi
1AKREaQZQ7TYktWS9LCDpTtpt4ko7w9NzfbjJ+cozll08pBAVS/JVWuuGEwdB6LM
3nZvSnA5rn7xYVFlkxOSgxyh2cfTmLqmUZ6w1vrnTwstZ0PaAPghqMC0gnfIFs9/
en+Mlh+ar2FY++KRF8JFgrNm3Q+OJ8YthfEOV+JLNc2vx3AiuR9h8/CcSOSh3t1J
VvC04RBej+D7WJdp6l21rxBM0W1ZlzEP47E3tSoq3YNGCse21t3KtlUoOxJjI+0r
L/5O5aI6UR4t+wP56NrY8K5zYg+40m7khtaiGjci0Av9rkoOgFlX8ZkSREZrOWfK
mFrvN5Jwy9sFP1MEO7I07jXQ+NB9ndbgeWWsFkgSI/SQrc0KfFAUU+OhNRLdy4+U
XtQkMPgMCnwo55kriGZwN/sCAnWYgSS/ijXPRLXg1C1ttcv0EFQ1FVMeablfumAw
E7xHkF0SjcAEwQDqgYD4Irmsigl7jqFG/Uie8A+YFzxUL5VIsYaeSeOp21rwDAYS
PTtUAvNU2idhlNYe2v182VfEUp3LJTqpw6t3sMVgde5iAOs9sl8sbQaWQlBSQPLa
CCMP2Bj9iJMBu4C69fRnNsF20JEvR3LUFcsgUGq/7AsHxJyX437B78Oa1AouFrVV
r+nekwNoavkhLGajsL4fvL2T4wu6HD0Uy+QYnZgDSx+vzmYvOXD407zmJ465QRYQ
Yyk+TZfKNUPJu5KpTG06w4rajlUlXrHXld5IHCIEfRvtSNRZI4oQr2MNrImCJ6qk
lKyHV6g5pEzJfz7v7GHZWrz33d3LFUHnqQookWPghw6vpLzTY9Is7rPu+9u8kKMc
sm7+gGc8ANB44BVeTV3tmvljQ0Y9hvO5RtkXi9mHkM+2GfW9M2l8ntgTTPstxh5F
HG+H7Nakad7BDEiMfTV+Cxcyj1QZl8O9SSEZ7ry2U6Cpijgu5FJF8tLNaFjEPL1Z
jUb94FhR+gwWuM8EGymGSUumloQyz7KxKNojJ8lZj9S0s0XZ+NKOA48cGJtg4fOg
psf/3eOpYhcsocbntfu71OCT/XzSZAdTr689W1HfYCcZjD0EHaGETfkYvHUtDlBk
N/NCjj19dgUd8Gsa0osOFFB6M/wWYbHsQlKrCmLZefViBJKpnd/ckxkwNK3nVnTN
QzMMKpHMhRCceFuxi6lMNJQdhR9cyGjW0GSMsodtuUEXO8rzzh7qowxzSOHM4sso
CgDWEiZbVCcKCN/0+TOSp59y59FwL9C5hmWBSv/kvb/mkXPC+juXNlgooPcI8yY7
6Y9RzG5F6lMM6O3sZvxC+KiuvA2tXQLZAn05z3d8PXIbV4/dUCnIBpamm8C6NH/s
AEYyidF8gbga3Vbw48oF2J5BCT0dR4zoGkStYcwWsLTz5HY4F1ocVTUrDh1DX8xs
m06JMBxdhkHR2v7AeeSuwlIoTgyRfXAgDK1kbNQ+KUaS+0siGldqX3a6uYSuRW5S
IEXM/mVFOuLHKVK/aWQVRSwCoAZnNP5nmhaYgrjRL/2fgVCduNmT83JE0BdV7cK1
hSOIjA3Qg0jkD0yL0sv0tDFgcMOlpeTBgFKSp/r5x4+4Ycwc86M2x+rMWcgLQ/PX
ke7mHvaOB1yuI1WOh33fFp6Z0AOEbOSXvGfl70kMK/yJaHbvHa4GNqvUGoHbuVT/
fENC0vWDxGZSeoV2v2aqa0+zUaCzcWd3wRszAGRC1YIF4ihpCqcgZiMMhKq193/b
ScdaDQ+la2PyeEfJ62+FKDYLn4qFrrdMY6hib/LVknhixqiQwe91U3fRoji5L0ME
0RaRgAFY6BdNl2aLjL/IY+SFbVBD73BuJKqXK9GIf+JN1PrFGebYr+6G0WdnxtAC
qcBFQYH9n6IcA2xgugFC45/4vtqoUdGxpD8ulUVaZl3XOqUVDtqCU0CFVIpgfE8X
6LYv6EcKH4t8BjmOqpZN/3tHd2nXWOvfznQAjueBOO3nlpDQ8V1X03pbJG+ebp06
IDu4CUlkqbvoj+kWvD6ViPauaYojlQyLjI8LTcXqJLEvEy2G06HRQSXO+qRhZyea
Ocyx+4BPisgDrIM73nAQe1NCrEANPZwKqkSJ7HxjRD0MPFsW6H2DUmavDsJAKe+Q
6yVCU9YqO3lcka2bkNUKvFG7vcikOWg19oa/PWSwcVeRvAidCV9fvV/qG2xrfCn0
80P+2FCF2guI8tMUvLMWMbH1YHdMXXCVHRb/eJIp3v/D37qKybIie//7Pb5IEWKj
LN+Fq22n2bLH3lpn7ju4ZDZu1HblZKjBM1NMbM6EEubHMtkJZl3dJrBFqB07RU5z
i7PGdrm+VdecLfuxlk1XbLwtDzFD23Stj/sBRd9FUZbbP806xH6eqt30pY070TE6
zLIqVqbG0DvnALzx6MnAjbmheUGRTRiK43bsBygJuNfhXW2cinN8YNxXlFUrwhpG
ZGpz+lyqIskzx+qA0mmDSNtvoTSR549XUCm5Ay9LlD6j4cf3UeSJPOc3S09d/QDf
c93emdS/+2cG4K26XiOXkRtY2ER5miffg4WGw5QDSGMrFIqZxykHTbl9BOWJKT7J
G9n3CHqikbCBSWLprnB4wBCVoePT7lOJ91SsRcjPq5jQ61SzEdSSsUdx+7q38mEk
lCp1Bb/vsXI9pMwDGlIDvYFV+vwxLDBktIm7XKto6NAv9NFUvENE+tBM57+8/FQS
XKtn6AqizPoUcMzVFDYm+ywAA7KQQAljV8TmzLzPTM5uFOo84VD98Oevq0uJXc+5
TUdsg6FfmdCjVaV2zYu3+uqiNYFxbSNWVzW2+iOjY6dtxNMBAdjsk4KptUmE7Qi4
wPdbFYt+5WJhaTFdY/Rs4Ums/PM4nsfviIUv5zVKeAyFPpRY1ImafS3oBBKsQ/gL
ZOtSV4BHbF8HHnC8dXMdwGHqbDXZIX3Lwdv9HGdYagy1m4o+X4dcuboJTqOuUFUI
iB04ILzC3bQ2Wmk/AVIGkIt4sr1u4JQZSeMt7QxtiOebJ7yqvSxkbT8RfFYU0lUM
GOx5D/yUI8sniFMtj+qL7ZtkOpRjlDvDQLxyUdE3GYysEq3fVdBfyXsaPaiO1sSv
PTqr47qOOrK8BKw5MSjc2vYeZ8FltdyLrROANoYUnD41f/58om2GZHvLgMTWi1PY
jcGh3fO4ONRUkY8U94s++G95kCbm090pGF7ssNiIilM5Whgcov5EF/XQbaeYoUGu
gjTh3MWlamuXEq/XLcb6n2ojf7kTe21f/wZ07wnuou+QtWLELOpexV/o7BOjIs3U
JqFuGC6KzsLOaz/w3OYrTseIpntFiNYZkn2wcfcfcgL+eTUlgwo36Ur+afh+smrr
ju9En+jOvy284AeZiofBzNNaNqh4kivVVv812yw1gllSLbHr3oNJfG2KdPQcYrSg
uVDbK0TdPoz+qE840zRr5VG+9Z7TpsvqAao1dcwVl9K1H9m5gM8Iuz2F2uV1EFf8
zwpw5JA3AqE56QcO2fBXO0PM75Kq30d6GE7PmdaJYDg74jIRppofCve3T9bprfmi
QhTCSAsob+RiZU4nOSXmGGOwraIFCF8jfn3weWDOvsPk+tFNMl+FsRIXt05jXVXD
RzzMM6Pmciu8lCf4K2y9ovm9MXeAoosNMo3V+ZNO9y1N6lxUI1+HkEy1hb2OXP09
NJd1iVrhwjVElUgpd8qDWVXA3dpiJLEXVqM2Bk1eC1hH/6rBehieMyuoCIhTlCls
uhv5/Ktbm7jYdazqoWFXuCYRYmYTlxLMps2GWF0DI9O9yxZwm585wf7kSk/vP5qd
1BbdXHeDV8T/A0t6s0n57Z4lrq8TXlIInYT+ngDmcsSPKL/qF4AvScR0UwhKLwR5
xGCgJnWZdfFlZd0R1ODr5TJ0QH+Hug7fJEGwLaU+ZzlcWG3R4jo4409to3Aavsdh
FaaFCgLCA540HT2TEJKk40ATUs4ym0Rov0tJ2dju9+MH/HFaMbwa+MLU6WOajcpI
8GNxYCZZ18cEBLAF9SdEhHpkU5m2WktcXkYFi59hkFl/ioCpva5Z267cQ8aXd02y
SETDMc1gAzFnq7RgkSVT+R8PEio49J3Uruq/yssQShKGU7EA5cX0TNjbTaP3EYMO
T/hFqnUgYrdUaAb5xDpeLspZ3jw/NlXCTdsIQvYEtqJ17jgYFIe8sNfibhrJHOzd
HmbpbmsLxJk3vZ3XaCglJ0SzVbb/rqheKdrKLaUtWoqvrgDHxCxhObMC89tazs/s
tRiqakP01HgD2SfIcQlGFIIusWf7QCR/KH2iveDeb0L1YM+VWSZJ02Ssz8+XR4SN
DwZ7MmZIC8V1IhOPmNOfoHebNT4v9pn55yV//TSDPI2P+/tjkj1qttAs+rZRjBWh
ANqZ1PjBGm4v1hAq/iSfJ3q5geN+UjjEqpSEOGOZhXWBd0J2euwLyoHy5H5/BhZZ
d+tC+pW3VtCeMrv7QL2wcrmabhuIwWahe87Ug9R3Z51/7F1KLlLzFHrU69SOsAg2
pFsZT3zgAdu+giMeVQjUg6GKAYblYSKtmvpSlheXIwyQ1f4do/y51jd5oHjcESN9
uWnAe1B+x8/+gP1SX8FseLC+/vHNMN3qeLv7Q/oM/rzXVreeK3MiO0Qeh1psLKio
wZQYlCM9D0DeexuTgpfnGiw/o9ytWvGvfQXTPRlyfUqMY5wMyi5t4bUZbJhfSOFu
A0zkQmUoZRLEI+edOPAlcQRalXDj/YR5SnYY64KNMD1/Z7+Eu+GzCzuopHAWLoeE
/hyop4rdj06t5FNv7+QqOKjKsdtCAndtlba+AfjeuYz+9+6ZbYbXQ5zt+oQ78RoP
ppYFECdmL8Ig5iSPP7GR3cu18ZxDemPlXMGwx0Mg4WfN/0crTNTb3VIzu4OK5lO2
9ew8d247tTsKDja7z+qRJGP7/75k9Qnk05UuHhOyt0ez/2S9nx1C+CjhlForxgLF
HM4yQMN0CNChyrd2VCIQTH7rD3TRw/1Ml+TunLVMQDCe0wZKZjJZnsscJcfjL22T
gotVsBA8RrDz+jG03fsTV1CdfAG7UFGKfvRGfiqmE8OAvrXdPBmiUHLwpM/Vyk2l
NHKIdOZp3MslqAxKKNbHr2lYEtJlqL4/OxZWQzeREYI6lx19kdX1QAAzEWDHoSTt
5BNKUUfzvIjSXRRvgXywHfQ/dzUAhu0aJm3Jkaa86GvdNnUkpDZrjHdRBd9jzHIU
heFHsRLcoDFkoLoojRYZVosvwlhK10fhsB0f6aXjbo7CDnxIgxvs4H+QIy/JCGEJ
8FiMgT/35GdVeeZgIhAkCyuSh9c8daJclLggMA6Mxz2cXcglb0PBEOsASCgSjW3h
R6LTZkgZ2sSUE5UlBvw80wwdvZ1WNKT+7ZOJFCQP7kBtHz2L1R91hPHSLlThKbVs
1RBhm3jinDfvWwG87HGwRDQJC19kCD7zI32HyG2d0ixqwRoeEtCKMVbC7gvPyLQV
Xw4/nM0MoUGIA062Gup0orYP0iXPmicqUKyNoM0jHK1sUMnt/t4LfE4KqCG0/DjO
pBiGatTh+XJT0iy+0lj8ueU44k4saDGZldaaFLbkCYs9iUk1rGhbiJmDseHVbZL8
lHKeXSZYTMHEmcHx8nKGSf2iKDr+4QvShVaw1UvlKxTXwuhzeBs7NKAGqVR9cksh
4+1m0cvrmxzYA8oModxNJKOOn37MOgrve1NoaNmrIo3wNMRc68XvND4izeGz4eyr
LBvBkFw6s6DeAual+tZvVCR+jURwI1QxgorRi0n/UoC8QzUK/+ik4r1klWkIgNOV
lArGP1/S9YqYgeKJkryiRRzOP+JYVFejnF6TCJv2qJnYIWK7zmpk5KQMH0jtIyEk
zkRF0J3FjjySKicS3vAepX0aJ1AvWklucUkOxju7ANBzt7YIVMOt1Bu0xy0i+/IS
eNZlKk352NC9c39n1ENMmwuBGVH3f9n9ydz+yqHVqxUpRCo0TZ0wuQkjCWo5LOT6
WpcLBwmk5H2afZ6z1HPlVH7bnx+RGNZdvtZznkQQ9OYj88H9fTl+No75tH2ZlY/F
h8REQKWiGQR2WAAwkECJcG+g+mjpIXrPyvi7vwtimAVKNGB7vBLxtdFo31mjfxau
+UT3aB4MZNVUwE3emNi9QJcQ3JT7tVp1uxbPNWHifHdJWSzBNtVoo51Qk0kFmCUp
C2Ihx3alCqrIQFOuv5U0CApBfftm56JPD4xK8xejOs51wLOtDSMFM67u/1836FGa
S1cYVshXoOpZoYdWHv6fTKUysLQtXLTqf+mPcG3u6Y2nNplTrp0xInpw8y9hBXi5
F82cNuPqdut3Bfv3fkakwB+AB4D0OdM9+IuEplyQEgUmIHXGmJTKu2nplh8WA2aE
Kd55RJfs1oqLsoytfpLLBEyOiwDvknFHZvHgOTuaROwxEejJlo2bslwWaa/e1zYR
8AMZe8nzwTFHIvAXwxHJYpEowJqxR+LaEfCw1WbG3L5VON38yRSyjSvnyyIU3RI3
5SbgKXlNbcC4Lb0EXJmhT9pceUf7Ahwum2yHJW3wS5zlqUAo3puQGxrjV4qjfKc7
29W6aE7kHpM3HjOHmHJ7+coPyDQyy2jYQ9/mcjZpj4ezIHyzPEaNfkrU4XnwLkAC
TNUpS70wzEOXK2Ype4tUIro9L7EuyNSzU5nplf+bS+g0euV0UEFG+VI2rA3Kj2ar
uDdm0JRC2uMzzt1nkhF7lxGIk5ouS0kMjbElNLnr1EytRc7uVsV0vlCxDIaQuLL5
53B0oSnPmk9sCEW6c6Yckhqy4IgrinyaNGZc2BwSlyPKZzpqci2tHLig0atmBKD2
yrwSqvB5vB6nR2CQJMG8GSexB5XVq8UjZ5kyBHVRgTAax5RGLB/vXPjk0zDMsXIi
V3+eQ4rayQwXpEuFTKwW7nGdTEUI86qhE/E6US66cFO80ir5PBtGKzDaGxGzi1oz
04I+ptAwdAJgQKoZsJmxO9kyM0l9OI97Ja11KC0rjuq4Cq3p767O6wQgTElSaBEG
mEAqZ26j5r6slaCLyXQrqnu+VTy4tdX+6tHubLgCBo+7a6OEPpR4UexlpHngahW/
ewShUjHB8wEvEcP3DLgCE775VDUwW7yRIGHs+ZquCY1pqbJMgQtZiEadFxlcFoPg
5yE9e2iePzsxh8/JbVCHgV6Dvzu1nWcR5x6S/8tKIqrXcySKXMZCjBOc00Ku0QJT
nzftPGMHVarbKNmBOGJEa5l0hdcBDxah8ANpAz+s8BavkBGNU/55QVtteclfGvRO
5f/pY9D3IhSuogYEqKNJaS/H5NyOdik5LqH/ZpIY5dCle4wWFLpUpOgFZfkmmPq0
zWuH0sOF32s+mets/L1z/saiXEHfkwmAWEPP+ogBPwNOl+kuEl1JFXo6a8ZaIbHi
CQHxOgbtu+FwP4f6pjZm7B2BsbQu08ueEiga99xrDmQG5Ad+OHEHkdWFgqg7swak
P3OP58roj5euNVbYtzuUHAmKU9+nOD1uuN371Gw4TO8g4qD6FrjaPmZ8SbsuWGUn
zpPcxhxUsW/Do7O4AmLiIFNuI3FFAs5fI6rvaw5aHoRxpEWjGMLl8sg2Q0/rnb1A
3F8AOyywmGSbUh8vsbrJvhFgWcpU+hQ2g1JtZwPwFafjGnajK+8ZZe7xOoPxUuRn
NT94/JDZHx5zru9bE/aju9DEyyyh9OSBOo2Kj1kS15p06KfIsaP6A9zrsZIpVWLQ
pTWfWGk22ohkZwnJ4O994YpqgbA54hRkeU5dDRp0fPHjbj31ayO2fpEBCzWF/IY3
ADr+uywBb3kGhS9Vizju0A1uKiufgPEykKEhX7MrLAfvje/V6iE6GkeXmfOtFiwz
feU5ECk1/V7jsUpgqU70mHB43crvoO2jL8zWpUBYfNQPn3rQcy71St5lZ+eCFpS2
Dr1J1VCSANUDwxvI83wa6dP88GYs1meHFeqzSbOMG35A7W4mrVuohdciJ0XZbFtS
5inLCu6w6MetFRHjRt90V/cim1rAX6TasJDaZqGOYD/Y61qW0LIzT3nwXXc1YSRG
F5XYYaTWfkn8ANDj4dRt3JINO7Uvyg7beRjz29Eo7OoXCPCORinDbTzdSxtYlQxN
Qi1y9Ml0P3bag72uHfedrO5QVIDewXzZK7glvz+a4Eo8VLtZHSHNHvdfWoacqo38
hpYkTbEZfSqN/rnrvZrWtGRxUcRDgtKg8VNTmOiZXJI9bsffNt4Sn5q1PtwM/Nzc
Xcg21IWgCt/6JaezlVY0hkyH8rtDiwrKAL4QCP1a64uK0qPyRZTK4Nuv+zuTZ49j
R92KZwQg3ndRO2S/HEG9HCbYeMnqKCRWmEfuzpdPEWI3namgZyiQlyzepIJfPVpC
rD3ZVX/pnS5lHRm5XEqFk2eC7zyNO8C9I+OgO/MflPLbu/mJ3Io66KU80L04Jc+0
Iey4B9ZdB+/q/V2K8qUZfPrDwRn51jie8cuBgGIUVYoO1w0/j4yhwjvr3W3i0Z5p
kYy1s+nityb7W/ON/zgXjQLrMXGbkUokHpItkYrYow8v2jEG58rcdl6fDf+rY85J
IzXUEC+Eb4ZmiILETUAb/y6VWAxo7QDW6W8BzfbydRizPnR4C9EFOVm+KdNReOAi
sE3J41Adxo5y9UFU9RM4rwh1/lzZx31A20OPfV/IQLNQDSKsZEFq5F+QaAbGMnBT
vJSGtXLD3IvXc6XQIEL0rWrlaSfxwfCaJYIyMRTS3qQbbKZAhlord+SIDSFSVluX
Ke2Ox7KZmsxRe+LW+AnScZwmG161yUNM5vLmNdVy13QrK4XwDkrJFkuVWyNZXOVw
xfDeVuQORAu3Zn8ZxqZRmVAYv/uo0SngW5KKjKeY8Q49so0Wa9I94ffSrPwGQhhZ
Bbpd4WATiRs353DrMr5vz3sbu0m0HgiuQXgrZn6ZggPWNiRoe2Pqi2nvo+tz6o3h
paf0Gix5VMTEU8EGIaYVIOfU5u98roce4UTdrWi4mNW8XzKzny65i0BCqEttDzxt
yWajAjLSRzm64CGmnYwi9jvIiTHThzK8yE630WCFQAfl47UhJ5GoUIjwRZBkqOJS
9vGyboXubSe0SU3rLM6ydLOi0Gtsqrjw5pwnxJlMMqhKSl+xMtiqDitBaLmX8FdC
4xbLUaPxMsxcxTCXQjYeYnnKLTfSbg5E1z54HZk/Trmxp50H33ryfjd/B1GGqXh1
O87Vbcwxa1U1sM5LrmLLghA4I53xuWoBiVvfLUdYOL1QUay8U9U+6snrmmjVqiY3
Emx0V2JuRVwtnNfG/b/imb9a0E//V+gBpqrETqZ4AIQnjipDLLMJRzPM1NcgtRFw
xcIj6YRlh7dbK+2RS8O1otnA2S6Q96o/G+sTDY57uvLQeUSjM06oy5YMC04rmMc5
gppSBBl7mhYmKbl7XUjXqvzETAHMpdFEoP93xeDiPAM3S6oh3IVrXq3HA7bSuUrs
VNbbxmGVr7T818dBNuVjnxqXGdPVa9gMMhqy3dRiDFcyQgvlKgmSvSCSi8zGDK4z
Hv0jRiMTABSt8dnyXLfY+ASx/qq6ujaJSJoIM8KLC0zLOUXrDWzD618A2kywSgdS
Bdl3nX8hYB+nYX304OmNOC5TttNj9qsXOiM5yshIGCTU+hys8KG0CrEDkw6ZVP37
lQ6UGx8J5WR2/33GK+ErvNc0e0U7xSPRbp6QCcmO+IEa2r5Ewlojg08o65u7+DkO
3ePnLO1IxZ/sYjA1/VlgqlEl3dSOeduz6RpDStPzko8dPXRN9BLwQjiWWF3A5NxM
VJm86YXOsr+fyOd21NDpg57IH/XHBwqC9/Qf2HgvG6US/Cf6MfvyMSLFpNpCaFpR
wrg72TyBfjZremsr0nbk61MuVlsKHI5PoUPMUM527KBU6060zZJ95KQ1CDy/cWYz
VTfzhv6yCpFOoIys82gRcIEXx77G7PMBaztwGNCdbt/UDuUSvOj/o23iWNaOBr5b
Vvq7TEDqpdnVEc0co8MPCcwRhQ7se7Z+8sNJYgVJW9kfT6g/hlNMT9+6cHMpOMxC
KM8L7hfGXszyTE+Fy3L75LuWmS5qg19gSPwEFUTw/IxCgbVNB/OlGMY+KGs42UIj
yUKn6i/J9hszISZRK+aFECnoCqKEYN4FI1MkNmU72lVlDOoNScTT3BEtNVG5Ac3Z
j6XAMbhlqpTZC1NTuk7hQrF0P2waz8G1wTqHNV2pF56dphT7tM7W0Duy7wLmV/6i
GmQEM+Kf2Y0vXz2urqHWtC6C7Rqv10otkxhnaBtFhNicv0/oKdwJ810UXGifHf8U
HSAu4KeAz1lop3Co7vLaacH7iMoMm9A57Q6KWw91pBCZ9+Y2ehDyPX7oQ5AUHOfm
HZwpTGA2nTWtE6Wwo3Ve63bQ7Go/gA9v1Z0bIGZu9qrjth61LUm2esJ9NRrcxEZn
d14pohgPx6qMplbgsRRPPWFNoDI4GYqHiNqGW4tdKsf3kv1Hg97H1wjy1REvUgEA
ZWM4Oa+OrHopHdjxdnmGbYvlUssXiiCrSJU74vgQvWvSoPp5QQuXv5i6R4VEBXjb
O/XP1JG2su5F13wXHV8FJp9qzISF+gBUO1uRVVjO3aKcja+uv5i4nNuYVCQAl5+q
/Ic3kFt3bPkDcpN3MUtXtO7K4qenT8TQy0RzVmY8fecGQJdCsDhpZDBXOoN+WKg4
zdPhKjBigmNcKFb0tas3kzE/K0tO/MxyFn7QxN9+PICQx2U1SPvWBOi/apkHGg9g
+tyYN9cMUiSBLTgNuHWCtG5Ui41fBSBkawgEu1E0Xk432Elyu7oxgyupIOx+Xh7i
Gu5WLVNg7GJqxEwvt/RY1sqk+9eptybfT+UZammMksUlUSECkbl5yLUll91+RNtK
m3F9TDVZqnK2IvKXhDcOVRfEiplXomVscW/j+JngWZUcQmUBuWQZY6e8aoAqfnTX
D5PlSJznXPtoRCwF2etLhGo833tZF5XDrghqa7qaewu07jbMQkbqrM34SgQUXwWA
podri3kkyxLNnQov31x9O5ztTwNzHfr+2JObEDXLH3QTSQeiwBGNhIiZADOVNzUr
F0KuwzjWD8opmS1kZ82uNWn0kww6+IuC7s7RcDDKSF9t/gnZ6E8oZi+eDRL0HYeH
65gFnIBz/cgvUXMrRcVcTxyhHfjIF+jviz0znm26Q9jdr15ppRO8eDPmL3ht26Uw
6/0BIWhj6m/6NvKdwoP10RXRFASnqWrbY2+jhTv08qpnpMC8jGTC6pcMMi+NV0Rg
FlAosOHmSecV49evqmucXWrT3ZfjD9fd1i/+yxUdvo/MyTGuJoYdy0E70/g3m+AZ
23dAQ4PUU4yxzKptAiglaMp0jK98Jjz6sQ68/EmQj2B2Dng8oT2wsjnxhzWD5pGD
/3J0rtsy15nSppv1MmkZbmXBniwetaZE3VcL7Tt7S6pUEpdDhYNrqRUPR3GlsUoF
6xJImslQQ8RVvQ4/HXJPkAKpBCfPYVxybrSTsrcJzcZMSmWPvkrr5L2iOrm/50YP
SckanXLjatbrbNWSbK6QhoyoBjjXsAPQV0tDJZfPY5G8CP7qQOyuMPZ3YxRBPllp
U/26UhsQomcEZnqGQy5VQu5IFc52di/go6Pxxwfan3+2qqkaXQVitFznJ8i69aJS
e+I0/0O0K3XCMnadJFvCuMV+Ps9ncMyMa+FXMi0C8Wxls6VzerYUHtlD6bI+8p2U
wIJyApmqEGFy8hYKGrN41f/CnTGSQ+BTNwpSPmC6uhKKwYlFsQXBnUz3qEjdd6IR
KnV9L6aT0PhMiAPoCQLZSkvYM9LJtqzeXQzQR3edw0R4STUQ3Okzxnxui7e254Ci
l4CUlbr/sETA5DDsMDyJsjRtmuYqC2FVYwttj637GfOJnOEqxoIpTwwQqa5Terom
11BIiemXf9VHZagR5fppl5a9dC68I8HsopPsI+c2Q2lJguNUYs0CfpgvPkAEtIgq
tMA2UCG2oKVRC6N+c4hq2qTFrISo0Kt/HINdSkH7nUOy+ZkVCEYmp9MT/fjbjpNl
+ez8aOJAVT6kn/yQE33mBMJYQ6lqFVZhmm6a1FLGaNLlSmyrRNWGjlcaAIdLAqSc
zBjrW3Mqzp3+FKPbb45K3nQlq0EPVp6LPqU4W82AF5cTxA5y5t/Pe1bxAfYU+ofU
/NbtrDd01Mpg5DWYdwOIv/bbxbjWEU28Lr8n0Nv1PHo1czJjIm53RQoxcvaC89j3
xLn4JjPLTxjU1oamk2aNtBgdYwYo2XQGexDeVP/+vmxSyNPpn9dM3qIDWEvbHq1b
Jl82b2azEbNM9S4KhQyKOAog4hg8LuknlaB1IRimME0dJQtGvV4Rsry3N2puUTID
zZeqD8BWtSjJHe0RBf8CFMY6XKgRiI550FZZsy/CpjmvDacIx0lRTet4UGAzt+46
qgbgOTsMYxzDxAGuEzfbJdXzaQDv1MtVQqM+IcssRH+/Z8wpxXNsuuVKx6qhtyhQ
dxuJWwjzF8UA5msEeuySi0CLI7XUsPu4hNQmQWMuP7gB2WWHR4D/+JhTumas5yB1
s1hsddxkiv+1PNNiQk++Rpr4kDeX+bXmkHE1bA7nAusXTgUG4zHUhgzf9I9LHALs
Hslw2758Ay7ieF+EexjzJzqtM/BeOlOXQ014/qysgL8mfzCResdLIVIjyC6JnIXf
b1RyIDqOdB7IY/JF0eS9+tJ4xxZalWHyQMK1Ppn3eECDu4z2ah8evqW+KSE7MbyY
6SdOulf23VDlZtvPJiyNK76gl1RNbS4E5Y/oFXAILjFmeX62G8hY891xdOXiQG/D
Yd8hjELCjoK4eAPQA2qfP2e0Mj/qEOTvxUgxs2LKzYjAhkXGecG663qGCm2+jetT
oHma66iDVcUma4l3tcJiedrwxmhda2TPTGAJSq1t2jvi84ZStUhbqTqLcwQnFINl
enS/h5hKlcSH5UqvqZ2i1PB3RO2+3ExWE70OR2Yjh14zdsiUxnhb8vJABu0xLU9F
MSz1q9neeNwPYskmFXIxJsoIJ1CB2+nz8eUi9Gk0l6ZOST15O2tNCS4nXKfQs+4q
juHDlJVfdHFwgtTVseTfy80eKF6yGMzP6v+niB1sXtQ0O0fFXYsEHuUuYPdyvo8u
ugYxMUVNYNNITQs1p995OzYFwCHRLBvfaGT42CA0QaAYqKyoSh1m1a4+tDt1xJuX
0sQfysEOJWkibOK/1sE32WXyKr8HP5c+ZQGLFVKlc+GQ2Y9iSCIsh8TU+R+UGC/K
lBQtbvnsQGqqQAod928EcTyk6IvSOu4bEP+jlVKgH3+k6DYU03nouF3/S2L413hc
4YfwxWclMH7w1A6cEwWgpQjDQ0XfIBNrwCUoiM0RX829/hKbxUTzG1sRQQnzYY85
YBLfEsQojI2WOH298Et/407n/AgyYDQnEBEXWDulJQwss3xajQiJTZSALutPOWkc
B08N2mn3+SMkzYAsLPSkptDvca2Ie1aefaPWT6acQ97HKXA0nxWmLI0G4r5QZBE7
wzzvGsz43ALp3vkX/lJHcKlkldbuRKd9Rpzwv/k72kI8XF/V1J/IU+EQ0lOL4Zt+
AjAp6JfLizuboPr1hKNvP2Gi86d8nqK4jgCu0uw6Ytq+uFUSGS2MdPVyGqar10D9
7YthQXA2YT++UmzcPPKx0Tx2PUntXLihzkAeyrn/x9vB2j0HFlxAJzg+osKHA1n2
P3ht2cHAUGXPFC083h3aV9E5WcEd70QITnbigkSMRGEiXWpZ57rtkXjR81I+NyQd
BKBoRKd3fwkiV26AMi9Qzn1wGAv4Gvb2U8kihF6r3f8bVX1h0bTbZGdRjClBdkEF
9aWWKKVFoYFylGTwIDeSozvd6KJ6b+uyGOaxkyVodlrGasKtQoJjr6EGJdBtqU0w
tN83s84vlXHtNLyVzmGU2v+tdTpEuu0VHuZDorzktP1b0ikaZMtJYMZbMVKiPg1V
4FUW0sqVkgUZn5P7Qfrc78hz4BcLnE1NG2Vh5ExW/h/mUwlIxTp5+Zpjv1CI+dh4
TWhGteyuFnm0fTOs/1BTxEflIFkI/wnRSynXMSEC/LMzUZ4hq8s08haR9e31uaHz
2zxyKT89N0niDlFM+H/pIylJop7fa8U5EfHrst4KyD/jFIouBx4DvbCFQ/VRFO5F
hr/6F8bD96FACXcVxr+juc0i2aH3vy1PlA0TB0tF7PJzbdpQfaJwEplw/ttcZul5
fb5tQRS/SgndvS+Oro06VY9geZ2dC8uNUIStmrDqfcXfjCJsA2RyA4jzH6AYFW1v
g1bALH5/IVuozvAGTpf1wYTQrusO3XNa2j9CMILhCu4xOIOa1CfgAW0djTfnKhiR
OUVF3uI6vjsM0N3G4SWq9QOIKyTi/F/iRBpZ61mhKnq2xmmqBG8+Q7J8Fz1P2IOQ
pam7DTehV/l17irZE3YH8eBUXmIH3agp/eqSIsrCkdz+dk3Oby3z98BvPJa2tGPn
045PgoNQStuoYprKajtGzHyi2lV5xJE/vn6J3pRh81LbX8UQOQPkrv2FktzHko2K
j2TYhlMwWXDMIwotn2gybtxp1JPBBqt6moXJeAY/N13j29vbOPDOvgpZBjFYj6bz
xBcOdKjouze/21GHWvkhc3U+HR9eWRjn96bSIhYoNtzznc89WjkQFHBJeeFa68no
/3aYYXkED7IF7TSH92bM7p24/O1gWpPP5C+Cal+WsKmQPq6XzuupzY/moHYWIJZF
ybuk6EMl+V/5vQXpvhyTEiXNqIJz8tAjEOxqQCHTIjAU2z/F3VhSI78zEHnUvDWR
ts+UBG5PwwHm2p59wRH0+3rtv/tt7353VylOWFum9VfFLIrtgSkADkxfRTUKmmxz
M/6cFatJFTWdeOVe+eawsfqXCii6QHcEuE/x0sdIpqHuhqlBmCGQFmNbLG2+p06r
7ybObhgCUPk89LSZl9AlEl1FRB121N9eWqMMQ+C5Pb7/vDXuz6ygJt4I0G0qUTLs
lQUDItMk+4X+27cA32IKRVpiQWZ0i4+REJVbGDlBH/tBULZEMZEPtxWhPqCIkzim
yfpy2wbLd2F3jRb7+dg/kAwPrBdZl5LuVOqFPGKjUW4T+Hm6oYe3L0okMMPPoCDF
3Gw8SYfGt4SVYvJ2dptCUeg3R5Cs6PdKS4cko11iKWI/1fcfyXswC7OgVWaykfLZ
IXrYejo6WwkzvNFpRV6Pxa6YEMuHGHUpVFv8+hM3meQZBeE7smQ4rcDdlGJmg1IA
C/NHVOu2z/RL61/kA9usoyyAsECIOca1vz9rviBRbJ4JVCS0MyKz1Vi9YDrwJDmi
eLSm5WM58qytQBFu1Our7o5kKRpOI88PWV5GfPgwZZ1iry44MWQdpr0+Z+ijTahw
lFeFDQunTmyfjqwNwkLYNQAQfHWA7H4zXLoSlk8JxHPmLIv2nNs+6jGZjR2K5xYh
i8mgA3OQWNiHCeZ3CfRa1YAkAvt9LXqgs5fQOy1ZNjB0bacAlzguhmKOwlRKBRgv
+dRGZ6tZcqMFyyhoV6AWMK9ELxL7JYeEVOvNlX4x7n3/cIKbmq1KFNXoG/uWCKJJ
UyvNpdD2nysrqUOt/5R5UMY8+BwuB/3N/NzzkZglYr3Lvmn3VAzvKGiAUQn4P0X/
e8U8TihfSzV1CIOgVclqs7aqu1+ehVObzu6g6mrdLMlGBwLROjo2nnOzyIefVcxz
Sp5x0gTZaijNchbXLqYFGb0ofX0/x7FKRmKhS4JNj3HY3IqkrxNvvxCSjLVvkqUU
VaN46VZdf1A7v23hTdpVimJjxDglQ3kfKpMSGF5Rynm163w8WdqxeVBOHIOJ69w9
6mAKn2vpiXCYgwN03rpFe7S+3LHung464I/OXZcGsq2y2p+CiZxDnz/suOMkkLYI
VV3s0ZYpL7HrZAgrGWDkDLlwsr0h9cFKtAvYPHEyhVU+ujl/ltOw56mMhjAF0vI3
bfo4r3Ok/MA5ta3haSpFmyUhLIs2oxwAUudFl0XCrqcSnXOrhVXkNUrqBg1vM6XB
tmlyFkw8P0TxFxQVn4n07ZTKqyankxzVg8IlWng+8CZEIUZS6ZpRwJMWRy1+04nm
nCWI8en3uwWHSQfrUH3A8xGOd2rSmXMCnABqW9O9Eu4tRGKL/rqKhT5pQzg+Qi4F
G1S6Kd8Pp17AQ6U3/g/5z9K/1PLXCP9qmFeyEN8caU+kAbjYYuWNZKFWFT1vWX44
ZGyXowXLweKH8xLUX/jYI8+bn2S419ygxOdJ4eRoOK5o/CLC2v70IuX6hBHHa5be
QpfekWsePAO9XEgQ8C0rBs29BfwwSUfiGZp+5X55qfFZpA8IGSRPSvgftF/ftPdl
na8ZCdr8A6oAynm2CIZMIaCwlfnMLFLFq+mAhTGBHG49gu887W1F+JF9qnOmsiQQ
Ac6Odq8RaKJhad+W+zL2O3j9NIc8rD1pO0GviUBMAOG9eHiysQ8O1ScV6NGY4LXb
v+KuIG0KVSLWasaamVBx0Dg3KAJ00gJ+dsPKxrkrQ5PH5r8IwAh3OsrPe1UUt7fL
UX/dl4/AUXRx6svmJ6rwtG6ykeoEIAsstC/yWLpp2lwvlYCyW4UNO0mvIz1zmxJ/
UHyEjWiah4aiuUctPn334YxIvha8+wMMMPa0G1BDFUSIegpO4jujI4WWRvjXgN9p
drggwes4+2H6VLK0ad2olQGZgFoBQe6lhY5GcSgaDtGaZ8pSpBSpKnMwI+HaBIA7
ztyAmMIyYvCNdqbq8Nd7m1ZzWu79lygAgk1dmu+D0O4YOnAJlrnGGu8iQC4ts3MF
sIXVELQpXpQWT6VDOOIxCtTqvn45xs1k332Ky1jE4Qy88fvUlud3ufrZmcbrKHhp
XIRIru+nJJcT14y0/e6sOW6OM3o1oL29U/VDhMmsudsmEkweWm0kyFyXBJO28Ocf
jgrmj+LTfEA+uS7yspdSmEmKRLXCFUQJXDTJU98gprxuaC8g9G3+tDz+5K/EXTIW
fvnq15laTnpWY7Pxt7Hiy8lZID8KvTC//RONBQDQsLZ5JFYlLY23sMr0CsXQ2kql
zqtHazXSmHnOn1Ui9fliC6LcfNveQcGqjlfdCEMcY7burde87+nclPh+GfW0lx3b
U9PDxCxtUIJX2ew46jjVgbYyZj91rNPc+Zkp3JEp4EyCiOfTjN+lApdvNbutxCyF
UoA/nhe7CMkqPhV/DN2MkdOEOExA7gWzXIvrfXYTAQjOFQwdkMWd3pldWQkKGG2H
iO15DX4v2QEEnpv9sHgIuaTGyzw5FLkX0gOR+xvmYEARztrKmfVyxWihW8AhPKt0
2qUDyqqI38CdTLNuuKC53OCzTsWw8qg++3UyBUwc1gsfjbs6JOHp4RYJNeyW2ZGe
EA1x7EpncMWDVV0y0nCqgDzqrReDaoNjuhqu5JBROfSG9GYzaJHOS5KTYtuzhd8v
U7gf8/8jeQDSJ+IvqHDbuMHH03Hz+MoG6aOS+OJwNlE6+CL6qUPKGp74BPB1yX20
zXO/npvm/KltiDuAw8fhhStNpOiRexQDKqIBR0XBRFML6b1urXEwJ5gqQDgRAO2u
HcRlqtwgb6Yv09pyLNVLMaf9xwvf009jUk9d1sfoOHOYLOv0i4VqNkxkUQIk1vD3
ysQ+nOEa3Ncg5huVjw5F4v55siR6Xi6/HhqrwvUbPoiuRvp6rzS95tWOFzMwl/4v
3K1Bq7b8+wjPmHB2qfKpJVulaYUXFK38Ht8pU4U3wYmErSSDXDpRR2VV0HBRJKpL
UC+AnL/fUmy4ypiC2uHm3ReQKchnrbDyhESXfkUA+lGZ3nuYQJOfgj1MX8QiYtM0
62tdSgSecZZKBgcZv424kmcek5UaktTV5YahQV37ZlhNAAbQz1qUCAiN6SKBuwfJ
/NqHWqEleBkYCBBh+mbNqaTFYeq+kH4F1TUmuYVrfN93vN/UaQsPH4kqa3AGn4Pc
vJLS3eMgcQMXzrV2WH1P94Qz+aowEiZu/lFpc159IGnxja62MauJpHVpOP12/W7i
4KLSrLkBMNd4b8XZedJcPuuiTfiIwcZpbHbfkXgMz/LUeUiJlOcy2/5ttVddzIXN
vP3qdSMBvjbuH0N1S4GRwcV9+mYwwWBJ6oXT3WKe7mSL3aPtj03BI4lsLAOGVzVd
ITBpZ+H985hTcK70hYOF0EDxR7f5ir0VRFuJkhkT5P3FtEvYdKPbvOTtLU2ZNVW1
OXQiqhaJ2rZ6x/tcOb0n15u3blmTJbRvdGPQryD7E3DOaziodpQa36Euq9zCffMk
l4Gy/GQs9k9ZKMFDNspL2iXHVf8R2amHRIimnyesoBB3lI/1hbB+38xOC/tF/0K7
P0G45HvFcNUriykT4xa+16qxtuojrYNtEHDHFI9/6o5GexjJ8qG44vjQ0D0m8X5h
xHWzuWyHwJhbDdYuifdoFoDr2JvWcnRPfi1S9xIaNOVJrZhIlMPgt0FcPVECwF0/
CP1LQz77KMBGJyOtbCGPCYBReom26G2iO62MYMw3aXr6X2Stz4f4zBDS17glHzlK
mTzLSR9Xxk+QS7ysnAhRaJXJJEEQyr15bw4G1XvHurXsMQhYZla1nkXd68UrX6lD
TOH65enHV+tOpo3qK17I3FV569CMG4umOdtV5rxbA+1CEnXlfFd4vmZ7YhIB4SdV
ZG4JFWeKavwNncqrzlnPdkbucYCAhZ0gwfJnjKvFVxZF0NQ7jn6iK4WQa2Ldvkel
KHSTmv7X1iW/yvjeVbWE5WSzzioG+yNyoh5f7d4iXDzTnWXE8R2jPgHuLYUKJZ7N
vmT1Ok+lzC/reX+JlfcsubqIGRZB9W3Grk3/1wnhrkVvXMZ1QvQALMdP2lUYz20W
h8UZMGtEV0P1u78JR5dbeAL3yYgQ1+h9tFz4RLDukQ3GyZlcKI6qdtcxROqK2TLl
rz0p3EzBwz9TwMuQ2gEg0sPvmmljrMBVI6ElVTFV+vQPMaCBBeNwe1YgASj81zK3
f1QecnfXPc2UnPr4lnCqMDthqPN4EVxoLmUL8LSRdAjhnCHLQL8wEYpUYJk6HDer
Eq5P162EnvOMScwA/AWo5s+XKm788hYx+3pLbHLCdp/iiNt5RQ1w7b8dbEIMbfps
P5/NuLKU6ZtR3lsDkTirsbvirQGBCToagYER0/e7kYkzceqiXG3Xu0Y7B+Dy8Mdq
yS8uWbCrdWsVEPAITLKxkwW6AFMwjGjQQOMUzN45I/Gi4RRYyW2eNbD/ZVlZTsYl
NB4eHuZrs5qb2y3Gx+rS2squ5SHEdNTbLL8HLo3mqZq+/+U/7FCVQDDn35uapy+o
IyVluq/9Jy6uPxoLwh7hiioaCQwFK9gvHYnJ2tFoNcwmAJcttfPofyhhlfWLhO5V
9iCULVyRuKcbjWq61SGA4IHzMaINaveZ7FkEfFcpbkaoyEe7hkqtW/6O2A7HyuU8
cfP+9z/BAjSyxry6j3Ow8JbCSJ0R45S9W4Wfqvl1nNHeHFhxnLfD1Je7rB5rrCUm
yx9ZMJDpLyMOYVHB7QpFLE5p116Ess3MPDIGwXj6sAkgn4s+kLeaC4Qqe2kgGsR3
piRmMNlldnGqRuH82xuUEIkA/0GTTPLdEgLItA8xz7Q0xkT5dNNCBQe5szNovh57
1kZqHc87FkeJVQBdj+gTdqMbrITGm+aD9sAKZuDxdxWzXGXCXg1/VPq56xpRJgIT
Seiv/jn0w7+Jfx/x+HB0lfLj3ZoJf20T1eCs0tdRssY3tInRTrgLm20tEOI42Q0S
0Q5hqcmYvcMleFvNPKedCYhJ4nQfSmV7QaXbE3wCqe97vcy8I8XhCwCOd8v9yevA
BA2zwO6BI5iUqGq4WirfVgfT6t07IO/8t9aEJ3dqva0MlYQRQeevUxK/Qrvuxgwn
XPBtEb9e5Sr07HT0BLYWLOn0wcQ6j74bfLRKmIhuAOEc5OogbVtXfLBtzzfOSaJZ
AGAm2rbKVsmk7RzdiS6TYHSJtmig1Mzn5+3gqCoUhwjYlXxHFOr3hxJIq5P1revE
PeOYNZFo5UyLxr+7kyeKtrr7wb9hxUoVEByUmRJsP9ycNkn36DBcau3Ah8o1httS
aOBId0ffmMrijteoGCucScH4ho2gOpTWgx0K3VWGXwG+P46Nr+j6jmLKDhUV0OFs
KhZ/XN/0FuAK+9TWpE6R8AEwVMOo+mjiKiO6m/AyUKBQnwNRm3+/I4qM4P1tD/qf
/DqZb5C8M7bvm9ZxqvniTntgyGC/c5hcHboYcgw0gS4m20qAQ6Uc/VxY+na5wcni
2sGQ4UTHjjKG9ysOgF26nQjSm20t9OGiZrtjcEs2t8MeagBKldGLU/KOF/ceMlJJ
HJpZlAci+A/vxYFzCngiEBrStKSodKHJBGlp3NS8xsuTb4ixYozLbjMKio60kMYg
Iou2pcAej76lSw1ga8ZcVBGUSZAeWF2u+qhaWWCu9ou6Vw420vbKGXtl1M13TvU7
CJx4WEkVgRADc1MCtS9bXwXuxBLGeWChHDA2FpocdjZGkuQetvoKIpStfqXaXXpq
m5mnq+Ewez0OjlOtUduFOx9hsADgbdxlDD7Zk8FArJ8Q52poXmMFzyJkBEHepJrQ
LYD3GUJ3GprPomQNbP9pnvVCEEZcD1FyYu1L1hQ/8hubIQ5lHBdwXfCCdwLqGkkU
7zy82x5tuKO1JSa/kagWySCbec4k/GRX0azBbprbPkP6CJdyhKa5FympOlMGLQww
DzWmd1Nk5+j9KBuFOy/eQDfS7b6Sl4BL/a54HMLFu1940vsaJ26VXLCw7S6dpbxP
wd70dCEzs0fVtTaOwt9PD7MfhziYFADi7ZPwO9ceUHYqV7LMDitIVV7r5wTIK3lj
an1lhRShlVesL88tqay0E0w45IcuYLj5jPuUmM5RI7iysrL5IieSzhSFSkfHqcqm
px8A6cg2i/vU9hor+icroMzU/5MdaInJfC+hFKC9IM5nv2MhpkSg3TQYITNq/V8M
8yer7mpruCg49YNBTzEC8KWeUtvOgwEcW8SO1wfWpC3V0zPQsCfzMXPD2NaB2QEs
40rwzvKLyTKqYZgcZaR634Cvb/ptSuxNG7EJgjoIYV70mqZ5ArTcBRA4xQnnFM/h
EE+8aeWquBnWS30fd904DtRuWVRwYCtmWzrqXAzUaYKrn/pp71OLRa1tuY+l8xCx
SC6raYT9qrdlg5EL11E2Ho8gMiGz69eDOC3gJiNERkkDd0bycthRnSF2YfD8NkeU
pPkpYKFgwEddf7rYTBTRj8tZB0GbVPhQhOF8/vvJJ9iYNiaP2PtbeplUcUiLvEQl
SgOzP8UE9obrTKm7iQLXAeC/VBWa1GB2iFLHL8+GLkDYMnP1bZ2oVs+LrReLe2Ht
0xAp9SBpietYReeTGvWL3IX8STaAmnuPiH1p8Zgeo1v2f7jKJy8HmhuIE7Auw1i+
jAy2T6VZ6MJ6iU2ii5GfOImZpEZjT+IQaPU+r+niDMh0R9Ktzn6UP/ZuL72CF4YF
FxngHo7HaqfrsOL1kNP/sINi3uvSA0PQcUU+ZbQBHAsgh2HjiIEv54nl1UpTiuBq
GzxJ2WYQ2N44wqiwHd4pTD7VPCg/+Hn+5TJhzo4cR+oJVTb0nOLqXcljD6E2+wat
IT5lzAInvJ5OEYcaRke9P/+tvOh+zRsDn5yob0ZlfczojGiTGyFbMP2GenYBikSH
URnbQQ6JhBtD08tMoABVG3S6iCKY4dobaVCrwqZKTPIdJsdR6licqe0uZApG5B/x
4CK8Wbf5ZYeApvZPUMwn2EnkexITKU30vsJ/vV3+h/B0uevGVwhqF418C10AQUOb
FwSXG1fcheJBzHHoUDCpxD/14Pd6QcD8RCakIA6Qk+YO9H0Z+QmFfrHldUoZeaMf
2q9zVKve2kIvn/+zffJ7OLdJVC0YyTrsQLFAgmNJX3XRTpZq/qA5Pm33sXz7M+xB
wAWL3Kt29kKhs/d/oZ/YxI4KRdlpYaZ0l9SAjRnV9SGeZpIr0MmaeTXjfIQy/dRD
CPBMLR8YI3981lMZXTbAKBW0j5C8Crjnv2oQ0sN9lEtJQtdYX8TC+iQa/Z/8/BzV
ebyUr3ZOXYAUezAwx+Hyw6wONvSIwX/XKUvchw9WHqQhcPXg5YCCAHDEZ+AKM60P
gZaRDuv4PGpQrgDMldLTjH9EQuvhrYbCMQPB5sbXJIRPU4WSkTRecz2CQyJgfQJi
6LzcoeRZ85ii6fZBr2yrshqq08eVna+Cmd34tRG2lgYdrSU+fYOIaW4f7/61vIbA
I+V6tSDxUyfNmziiBYi/T8qO/ZtuKnS+6U8eO0mnA0ea7fb1JIDrM0HMfUqAwwiQ
++flqffmJ8Z/GrbDeCXBZ60dyIMlonxzf9DUEYy5lxEwdUspJD6oel+Hxzi4aE8G
aNFGC6wanASkRTjwe6lbOFLoZQ3JoKcQOQStRFZ6uDEDn1yVTJqdVj4U9U8e7yVC
aSOP4QvlpIBzyoqWYAt+ivKWgCATuWaL1RPN+kzfvcqR60ztlRUe9cU8tdBVwQy/
hnFYY3l8quRdLrCDDvoACP+eHALBO2wJp2umAumQ6kgpbqLI9Hr3MsaY2O5+m0h5
Yt5Kmy5EFBWYJ2fuC1bKQeUcagCN45ypgLqbHpuIcFZtaK6MJOYEkezUcQBbYVNY
2ele2TmrZttJDtDOBkIlsnfVdX4IgOXIlXwVuJhBBJ7z68J3j0YECiKbBd9chWKG
H1S2INn9J9r8ntSE2cjuWRRRgNeUeq5zH9xtJHXs9SMwPil7mmV5kFQxJgeasYib
iwQ2xaGbQ/xJaKoXCFQlDceni5DFXIkUApMdzAmJoS510Py6EiamBXqU0434DeZK
Co4uI0l+hhEK21+PBqmNXFZilXTzdIotGlHl83l3nrr1lpQ9+U+yS5Lpc5rnpLbO
nuGeFXa2VaUmiIoyJXhyuz63jZp7LgyxKiDuTupXS2LHYlIdniK6rxPnh7tVBtj9
vwVhazLte56UprhrjK8kSOaxas6nvSHqo01JB9C7Owpgpv2Ir0+yHKKFAGUX6qgA
Zpgrn29fs30LT3FXNpUdfxU8ec7YuOK3rIHXkZobdV6BKhcO/9QuqkEKo9a6+Wiw
X6lRwk4BhXAlEK+axAgRuQfiTkTBS97+UwzVQ6U2asuCQxXONyrINRCpwri0XNp9
4EO/1oBHWK2i3/MhmdLw2yj1nC7anF/Oi0qJ4UopQt1Fu0UlFq8yQFfBDzTwu/GI
bLF2sHTY5eBJN0Jaix/kbvy9/BMi72MVPClVjfPsKT3gXiw7k6JYHYycNdCDuUVl
gs0kaUK0KZzFpu0mz7zwJiGGMoM6SmtazJ6dvkBl2CWEtwChYYC4G+eNQKujuPTM
DFzhJ9O7uzpX1TURB8JXG0vDafCGMnoq6/mf5KMwtEMO9zsJh+/a7HBR+ad0dwiR
YPGDzDdYg/I+K3a9VuhBeRbp7pd97cMrGr1/MwWATHe3CGaxomsVWjTJ5UXBLFwM
9Ft4IYO+zAGnFeQuAgAn+rdfScMQHExyZY6fm/47jsRxWiwciEEiv56+s01O19Iv
aEuln0lAvpMSEsgOUn/4o0qTCx3RTlzLV9Ab622+KBnWrmh4M2B+OoM49BA4OJnl
2bk17hjlXcvjBkD98+5OBOHExYp54Tm6UxDVKtiX30g9zIC8v8wD7Uzp3uxy/u5S
wrudx2LoQJn9X5fbyxEUWU0lP/ipPwj7p+Lei2VYaJvporQnhugERCIX6yKemcdP
W/h/YCjNG30rUNFVO4oer9QvFdd2ua9Wp0K9Wzc/y9t5k71wkWrl0/EQmfVB7dCi
qIETc4W3nZPlAc6JygcchgrZ4VYxhV82rpWiKhm3kuDKYrMFD6/nlhifyg4+zW1e
yaseeJYJ9Rxi6ZeVCVvRKRXdQtKHLf3fFdCrEvCYch95vivD7A1FU8t2EMbfq4Yl
xZZIZxdrGg6Dx8Kb66/GC9nL5HVjiZ+HMAvtP9XniP/Tir2qhYtA9QawITPn8+3R
kuShyXij7kFmOb+zthCr2GA+IoYq78a/QPFjCQVo2bmZy0cEq8mMizYIgptTWaaB
aeI6KQ6WPu34TvkjX8tmuJa7DOPt1stmUqnGO2TnZuZs62ACKcc8LVE+K7YEZbDD
01Gwri/UyqCjQkFlJ/xnZxpq12uqM9tixox2LHs3wc0fjQcogZjSr+68ohlwHac7
ichRzPJraH0HJwe6mK1K/A/zkundNmzIAWCeRQBslu/CAl6YPk25rCHRe8CLZzQz
alO55WP5njlj4x6P1b5LuBnJaN434Taa6T5rNDugYdFGyNw++VXUaFPmhG7wFWTk
UwDRWlYLRxC66wneEcxnp90/Zqaan61fk474WKu2qxPVvf+pDjttNkB482cJOYcz
ooOUKV0YX3Gd8i4GMaxtioe7VPe4NC/1R4V5fZfX0qRHi83SfjFwbGeZ6wHrZHAW
2ikEolKLHtsAGSdslBkj+gCQJWdHzL3DKB9LVq5Mq/K0d8Qvdr5sCm40YIPYBbYm
tGintDyOKXozq0sYNv1PXqwIK2Rwb4wiE/ry+OepbCjagrA/dGelpLRdzmruGsAi
RdGu/aO+lJVBqdJ7WbbX0cvTljxmv/S8QWiSi9i8wI/egJh6dEjn23yznFLD9moV
f+C0rmSH7ahh6GxnMRdWSbI/2U2mXmUndYsJWZq5JcS69S5JqAzp2QhQhw4Ofef/
EpFkEdRaTKfrJ/9l2zoWpzw82C9f62oaBUZ9AFfJtdPzqhS0MUs/rXi/ayaQRl2B
FVjvLAoJ1yob+VLEfikA6DeOCWgyP+B9QJcv5IrPGyrrOON8cfUPS5ehvFgpQmRS
mz8+ociMR9ZfPwT8PyKQBDdsGBGCVu9+K2JfTSRLSpPSme48Zc6+U9MGyrS6EJoy
kd5qG/uRDtF0yXYLcHStdPq+AKhplpIOMrxMbeygbf/QgkyLtM1dteTVpZBfscny
+ZlEKEfpTtIWPzc92yUPhTuPJdCPNPjiS44uO+XNtv5dqSNo9xXcv2re8awkiJaz
8xQOu55y2QH4NLOs9Zvnt/a6DNumYneQ4hZkpD3bOpfgLoEnhyoRoNHYfklXm+IS
wpDQqKPIuUMmIzyrG2h23qJOJv7yOGzOIygG0lqj2Alq9Yt6n60ygdMoZkwxdSUZ
gEJnkKxmubPdp9+Nuaa7hX8Gk9GRFd8mi9jW8IiySAwwCkjxxRppxF+9hH9vB3PU
r537sF9XA52tMh957TtBNg3g6vrvy1lc96OK1uaZZImUvmSdVwo9kVSM4SRW5TcW
DpQKY2h5C4cMB5rdCV0ga4gURyfhmMuLQvEbVnvVaoL0aI/Ibd/cqOZarnQRFZXi
G9Ulh0oIcBtlEtzBoK7wo7hGAjMTqcTi8PPOcJHLfZKl6j4TbsrfdTbpRWEQeDkQ
Fl7tr6QZsbgjcnMD4uEuOkHb6yqjXpk0KZByESTAlIFvo7hEaED4IVsmSnmvChMn
8PuqZf8wm94DV4hxUSOs0hkvACYh5TUX8NT/urVXENGxiXdAEoyAWEy9ULW35jRb
1tRlwUZaxJLs5L9b015h8YtVry7emhQQAJK6HuXXcJ7zrcMhTZ+7iE0vidTbojFx
1MvmDgpQJku16utdcGXglcrsvCSJEybRgM/j0pKQCw9Zg+qOgo42Fm+fOOh1Jpc8
SmQ4TuqR60sci0DCzhqZsLUBSGExtIcdKRZn/aBVWFONCP5s85+XMTQ9aVO/Q1rF
G6D08StkIEG5uFRebdG7FZpF52WJuK/m2T7whwGNYPTGjIBeoh7DgVaIh2k6p4/o
8QyTjzpShikR5P49eU0CpLNpyCraECJxG5+a2rrQpXUjm5WNHlD4qPUqFSHczDhG
YvcKdSUmi9v71l8wDOXXxJeRMiOklFvng/o/uCSvLLCJhAR6Amt2G7cQaTTyarfq
VcsrXSAdPbtMszavbJVjTTCNn3HV7iNXwsZrs7ake4p4BRazZh9fxqVhxwzgFARH
xOR0AGFjZaGzDsPxRfbjkqCrHLfKLEbo2G4hu5ruI8qEHSldjhr6PQBm6CNkobmY
nMBVW21/tEUA+HET0Qa3pWXMr19D+aIaStkGZzlQVSCMoCGhs/cgQ4KwOS2YHNFJ
NTOdQZRRpxs8AknEjwM7ZgxArnMrvf7+esqYsrkIA2QLZ5EX6sAOjQt8dZ+zyXyc
batBtrKZH91SOMcO6fyBpZW/M4d6f7lUppfX8ct5rJgZ9w5sWmkGUXmO4vSC56Fi
MXpI/9inzycZas8hc9s+saNweYm61I79E3zaK8v+r7kcpHUm3D5ZQclDFCNynQkM
RaXBuVrecEM+6R0Ff7mBDxwT/LJkU5WP3L+DndWnY1Fu/XoB+NHjG1Sn46ok+zam
FRTbnIyKKj+3QdIkEIQLDtXpGr+xPqTxvg4Lxd8ePyY+wVVjNZrOTqLX1KVZ7GMV
KaMiXqfh/glu4CADdTR+YylvuVSmImIk7yeFAPO5X7dnYSKhETv/TIhQ4SeNrEk+
nGl4lXrKYVry+gPHI+c9iexeXL/B8RunyG8V4Wu7u8tG8EysUT0f04VXGkHRbq3m
ofvCkoxLSeO+YUnflvtiQpK8qUHagfprTY+bQo/xGi8rqRoE+niDSakU1dMxyKCU
TniU+eJnEBySMrMNpSK80r8zU+4xXw7l/rqmuPkioEzpC7/Bu6Hh1LDY5vK6YnGE
mIvRncV5iGhsTGvB9URoXocRkKCn1GBEXpHqjIIfTIHOOevN5GY+6znPjw5CTwrn
uzogm92ANk6g4utQ44TF9XT8mnPI1BCPaeoM79+i9u4dnAnh3r+t2S7bvb0dKjla
cLGO3w2tMdxALyfyuZfDvkunIa4U+Zwc+9jb9WYwwQwTbAz6xhZJj0WX0PbpbjSB
v2awMtsdR3riQqVZjqr14F+zEuAQ1QYM5YwHYqPvTBQL9/mrWtLXvP4K2H02Cpb5
OBK61L7/PjOYop8qGWjnN+LqzJkrYi7uVi0WeSSlYGUNalCI98Ey1sf6+tysOJBi
nL+Jzln/4y+JbuDh59QAM7e+WsdmxZaYftMk4q3rn1LLfVMQht32FgUn6xleXoTh
MbYsLEdu69M9LsFOutXIeeBf9DZH+iEAuX3vUJjYyBpO05o/3S8SlYBnFJ4HbM8F
lY40m2k9pMRr1v2fPzAidf1khuk4uk6RC1vUXDnWus+2nklnd5HG25ETCt33yQjb
l3Kh+fd+h1guBHyywiVAEltK7pAjvRDY3/V3YTpoSVjlyQyhdUWsLD8DVE1MT95J
6V5QOwDbUcLyjrpmaiKofIv/poG4DZ3GSO0r4Q8JzGkRV8d2my7LJE7qYUcRnbef
F9kZ0E11yYEyx1VNWlR4ST8aMU2YnFUQ1dqQXJjx78j70PoObEWJotEsMHxOWhdn
m9Wrynpz+FWTEFsnMlD1TSz9OHuWil1QtQ4l4eJa0bbaRaRUH5/c0KMb0Eo9rm7D
M5cGelpvdGUswlRzKr2/yBEfaL18Q7z/LBg16czYTD+i65WHMIiPmjhXmd68Imna
NqrP2EHqdaNQLw5DFNf3r+0GDeSqKL0jKh1C9UoQXS4tMHohjeuJwuGkAFhLAHf1
x24zy1Dzjkd1SDbf+fAeRdrzk1s6WUjnxfu8GgE/nTdwN72stJwmDzpzSLUS9jwg
RYmtfoK3CSwcDlcJFV6+4FF0l4XLK7v08ugY80bUUkzlC4T8cFv37C6T6ym+hgWc
ef8RxVOo8fhIzy2aniCXQ+hKfPtpW3A6OhvsfD0INODRGr1oGIUmxJCIbpgHzHxj
47C/0h2YdcOxsnUMwCy/Obm0rLTZ/pvRGSp9vytXeFrp2/EIMIWYfH/WMbs/D012
P2K8TInHA97acg+i0D3q8HBmGw5BKA6uymHDMaViuITQzQ9rEFgRaj3WDVY6f1dd
4Yfan+INTp3aah5vTVfcFKgaO7rcIYkglGMUA0VNp0qk13EB+Y6spf/pHdQeD/ta
qNsX1758XT1BEGEPliZ89+Rvl1NydJ2fHQml/duHypY6Y4k7+MDpsOvjTk5FfwMk
RdjkA6P0l1SoQl8mkf7VAtQ3TyuPHIzheo8Sri2V6VUUbH/aqTS5quHRzytnds78
W/yfkezIU6BAVbbus1+/FPM25EADa7vzs12+VuBbwoqLkKrAU1OSI/zBS1C8vccd
QoJCqWAnb09sTfV89k7Vv++fp6XgsVNn6yu0Y5kzGCUGqZsORqYmU+de9TdqnMoI
gDzvZSXBhYmhGJ21bUUMQXQd5wyi5GCUrNNd+t5FfyZjbXG/h8ZIBM4veAvO29j7
S/ARA2Qgpe6YcWa1E6dPuuuUOzOG71GOhTx3YZBgBWClVCISFQ434HgyhzeiGO3S
MeTxEJsgB3oAqdAhv3Cvsxmt7okk7n4y/O5kCVTGoiQeTIlIEjJRR/Do//JVEVcn
+sWM0CrJfyIPcM5KxPnuA7Cgo4TWNeC5SVsLW1lmiQPLXpQr/P5IbFjsO8UmoqI5
McEVN7JHKKSXVvKpQRCgUWOAKXwgTKAIAPmW70+kNjTl3vqOT3xCd+02zFu2j9Mx
lPX+KIOyqhKyvp2lwYUna0SvJNnVw0yGELRmhjUZrmW6oyLfPzSTiQpoimhHnC5R
kz5t2m23WDNtDkn/LB4wBVWWy9MkIyKVWH7+0Cjfnl6i3EC89UgMO5AHrq11ClwV
L4/iphffVzCzhH1qBmFAvbK9vvfbjRQvWxk8zXNEnEDgkq2CzgqCKv624MEDeTdw
34vc6YgTuynqFiP6W5WQPLmBXxiUStjvIxIgrNUt2A/g70EqE4tlslv2ERYWCaiV
dhfqy74c0yJ27GVR02A7p7GVGyd5DIFgk/TG6rokCKxembyrXxCYw19ynRzvAlGh
4wyFuV8e7HwlbcyF3SQnC0laGI9R5QPYBbo/QCeLAgRL3Fm6uAlOGfSsW4oAptzy
CIEQe2nK2Y9cU/YmFkadmyF1QLAVAdPZY7RvcJqXmoFqkt7sprXIKpgYPDPsaIaT
/N4Tjq0BWihbX1qywzcRNYp0PXcb+RrQHSrfjzRonyjR4lb13qrLZOo+sM0l3bBI
KIDf0n3c2HyVLcLTOfdmdhPKpmMemgAtqipAwpBEUvh/YRaVHd5wUr/ANRR1aXbZ
dF+N/992BFBEdlPO2/cnOCx9tzK5K/Ew5+8Eybmu0Qjk7OhRAO8V0/mMtasK60Lq
BbfA/RR+gc2B50ygk62aPVp3k8OGYnY/sqYFwQ2ZoAH7Ne7K4WVign6hg8sUZFA3
XiM3B7j8Jhl/Fey9BdPBj/X7NVYc3xV9Uh+pi8rAN88ClCfDnymjAjA9EQaj5bEA
+5mcp+BuwGixSvyyOvXhnGhiZysLCf9WAsKE7PaT0uTgoZg5QAr7jWuKLUy304j/
9t07VgDr5Cg41nfQsmt2P+pAXG//mSuYeI62eaYX2vF4QNJjGxmfvPn9vDzQHCc8
H47UklQqgw2LVccps4WTMjd5h1wY0KcC2ym79HSxmUFDA5CjIBE4Py5SIKft6co0
35DHKQVFTJc31QcAan12waSxjxZBkGr7+JHQTu/QDrkFQXCJmf5Q5whfylwF3o+8
1QpSFrX7qXjnZlJYDV1QWZ571hO1LmYW73C5lJNt4ox+xVVraE8Yqx4xTaGDQO8d
opk2MLeponWCnNwoS10ew76HgHYpM3ZrSY9dNfCo5z3Sz4UUkI+KNYKJz5eZkLW3
qvdpxnjjLmFO88twWwSEHWgeGh3gTAg2mfvE+HqdkKImgjliUVK97qXzjb9VsFwp
neFfb+tviWwEs6OYbedAEDw1FU7VqiSti4GMoQM/GFvOIsSgSlsKc2zp6aG9QpHG
EP+HRUAGfG1soSh4wUWETqMn4Y3fk0EzvX8cjTPs/+TP0YuRapwXuvgauOnvVynI
3MaRMpvFfhDHcuWwSPjh1TjIaNuSQ+jIUigQBMet8qq/q6lgnbh5Gfew29oprBcT
7IAJcCm72t7gcguyrxudXoVeyWynQYg9913RqFABhKTb9OHzhLz0sZ/JNlWuIx/W
8Go19M7f0AInqgnlxDBnnNv55dqKe6k93v8/UeMZGhSbKSmbU216+jnqHLrV/zWd
d7nKYhZukGLBcYWF6hrSV4nCtN5dcBzbgRGgrY8IBa8UtqbHFWceUlesATNHcPdS
uClchKEcbuFEyPN0Klt3pIwoBiGEWKUTG4owDFBn8tWbYX5rfeZNvFFYNWt29cyi
4W+v9CAT1MeYuO7bO06rCuPasqpfy1e/0R1nwYvY/QQeTb3SpJwKsegg9vjNYH3I
vXEjSXVTo2WE6IRZVAzX9u0kBcWHicIW9Kkp5GMrYCre0tMTi7DSZaVr4Fcy8b+T
84Uf6jaCADFSD8Hl4htHGN64cEkKaFB2NOsiGerlsKYdzXNDQopv6d5CsjL94RBZ
kuX4j7/ABJchMP3h35OdgKtb30wODKpESsUvdCfmRuhNgGkih5QyaRVcnHLPYkT8
UPy/V6zeUMcWqB+APoTFvhT16zkGC/i7dXDuc9xyvyzueni0kllAqBtI2BA5N6JC
NCfZKyDgMoEglmaShne9MHxZ2e2L8vUFd6iiG+u34yjkWcdTEvAnXQQwjQdLIGY4
5Lvi3U4TfRYKJK+LWlrARQAr96dOkMC3QQBv50C++rZgkuQX8AQKsdvJFpcwrg2L
dFlsveH5n/xpxRkj2iguSGS/1hp716nT44/MsGlPU5LmOUdtmXJDIj2t/CFmi/Tc
78DZdCEpbMA4gry1o+WUNBfUn1bsMfAAZOEB9cOypCtlw18/zehD+W959dZmHt1E
5lLUGYqdvv3EtGXuFhzuGm/lCDc2qgLGm97j4wFcfpNmzPsAXWNmpFHVoRuVFfcP
CHpGCQO332ka8hvpsLEiDG02S4N2APmWrMqHC2IaLorrpQ8hJ6Ktj8RBnC1NoZo4
909zMEGDyLRdTNThNrjrT9e9oZ/McGHeRYp+lwKLAaLl7mJTVbHfT1ui8XkA3Ywx
S5Y7IvCMIhEeOgyOe1E7hrvmQBqOX2XqQJsTXr/Nkjp8uHNJrz8NDzQzJbUFKy5B
lAeHRp+jhdg6J0vTe7PlZbcOJhpBtorG0MOUCiafguc3X0brBUf3aHdKdFWjeATY
jKetWQHRHEEobooDNFe8oCK5uZ9W3QYV2JL6Fpk53ebpbRfKb0040YF4wgk49UJI
gu93/C9qmr9+0MBrpDUbOkvHtaRmfkmynYf6jABIPCb+f8u4+IsjaFddGtxzrWed
87ikhEahZABK7df75vKMmxXYdr04P3iBYTwE1SaGCjBaAb4qYXnI7uhpED6B0/I6
UQ1LZeQwufUgH6it25+TckMYbUfHxi1JJyai1nSr7ryJH/cXRzW0UtHhEWbA75LM
MJyiYTm96yfbAUaBFNXwKXCmQ0FhanZ9580zUE21r13g7CTM7bj7Q3W8Fa/MX0Yo
Zi5STNiUO8c0oDUfecu1S+hFs7kAWywTKa8Wh5KWddKbe6HI3OcGgKtgIBOpgjMv
7hp9xeG8W7solyO0sPFEcZKL4NxQSDMA/rkZzRAJK37WgmZNOCw2qaKrOVyzOp5d
l832Sn20ZsT0ROKviAHnCoJKO3Jll27X6bC91/1nrsl1bJGUklJKVd1XMxdTizig
Xxopwji9b3qu3ukkwOhLwWbJRC6p1+IFApHWnlaMX8grJtXnc7TuXIDvr4QFTTCh
YOx6Td6bbFkrtm0ZbLyq31ZgTbDCxltHJOhndiFV1DBlt49prtyzm9dbd80oSfg/
7+QwsB4ATZThnI3SPLABbrhc+jawZ8LgK+CiTcWkuoLACiUc7h2m3XHxEx9a62z0
uBTyj7iA5UZe8ctNB/ZqG/IgDIc22JDV+maJtIpk02aagkyzQfsK7Oo7LbC8CnC0
uUEbKjqA3ipyuGivI+CCLt80d4r1Sn6za6p8c5XHDSAydqDYKHcNZAN+lLbxorrN
SAPi1//mbL6XnILFiV5bHbRMqY3Cdc8XzOmeQ2dxbHTZ7TM+IU3TDMOnjlTajvPo
wOVb2pHrmbJEEINqnYC4/YVtMyl5gs3H86tN4CE/SaDCZw0hHAeilxyMbuvP+awk
7wn4IQurb8vR/ejAa/TB5OqDk8AFDdMgByVwbd9e89AySaIb/hXqyrXcWrfC+QVM
CXeVWVX5y5RjaRWJIr0bAdjUxn0oCiM6sDK2UWHcOBN70hpGKajA1k/w0g90wJBN
24L60EK95VyX0SDZueKoes86EkdVCpJ3ag99z0whTc5/pHdTy00hIvNH/MT5DrGw
+yUAq3ctndHJGl7lR3w45X6xL1bhV6mUmwgKpUOkM66yVFY2KF/na1KI/cCj8F/4
QNIBor7+tLd6/ioElhenSrKFspGhgw4OtULKzl1LMxI2biMlBm0uwZEwmsRS7R9E
O6KJ1dIW2A+y8G02/B2QubeaRAX2eWMZnPHsTf5LLbLEOp8mxslWYzobx8LNlEIr
Zz3NRMB4V8icdFf+v2UDF+bIGzsY8Jg4O0jIhxyAyVXpdY0WVBVTzpU1yiH7i/8d
I0kSlcMdGM2hPST4qK2MYA66aHDkFL39IV0USJTrvQmxWuk1JhOh0j7kB/To3q5X
uMXBsSLKYTwGr58JLolJjOw7bZf41wfaP+SMvX+M/m8jrHRgmbwI9Lw6MLdKuTgJ
iWK+Aprh4ZXvDPqsD3dDJCpfPThB5Wjt0IjGLfJq8Ssv9bzJr4wk3L9J1MtH5oXF
0p/9G67smrfDBxue1bBkvr+1p4MZ0ystotgc5PLkBtM00aoFkZFnEoRU8Mup6HTU
qn+uHmTa/XMdNRSBQA8oZM6/nbTw47NMazquK8OK0QcHRT/MYomnl/5+cdUCzu/v
sCb1jIDBqsiC69iIN5EB0WDsYhxT8WQurp23bBWv/sVlbDfdL0rgxPgWAfwhh3Ii
eDhlWVmLUcNuWVrTGMlFv1VizeABkF9i7eQWJ1le3UWvQVpvIVzxdwFTaxoplaGn
JUe+XCYriiMPcEQTD8pV9GaEkb5P9EQ9LO4ppACE+hmEe8L2zbjfll2YPCEt7rpO
+qdYAJAfwNL45d/8VYwuFkbyzb4vdnk7mpwcX/hY5jyTtRwyRSCGXBQGtnNLu+SS
OO1uWwRzEFLfG+JoTCbduuafzE+W3m31DMeymfe3O/0azcrUmYpzPPa9CB2qeFNK
VCspVIoYz2JtAK8g6Bkzz2P3JUa2uG9mcEY1Ugk0fPsA2WorepzFOkxixynHsRZG
+id3IW8HM7UVL9YF/1vJwRjz51kVDbbncwfJUs7FJDBw/J6j834r2YSV09XdzQoN
EdbAMbL6f3A2OMjAmS/lyioCuBuG/UPcRh7j9jwsH7h3oTgn5gARnzOKrKnDJvTu
TFHIWm4+WnVZ0qaS8ut6hQfIAikE0CbRp5i7NKuYsr3VfxhqTVVuTwqcmik7+mIa
V3+qFoPpUelNmE0sPxg/3wk7d0dt9p6b9uuxaDsDW03q67HD+/+NPg7qdGrOqhJ7
nBXVKj+RkT3RYyyoZGBnswqH7MgnaekZe5JzVfwGmwJXTw+WxFjH0kz5Ww9FWn76
mLJbn4Y/d4gCw6YwzNuqJLKoZLNWiPiP1EubAbsEmXbeHdVvkOQvnXaMyTEJ9rEM
Ml9NbgivvbrmgxVnWTOF9NCwjFlbhakeLltb2Pz5RVSn3U6m/iAahRyE/muHSMbp
wt8P0buxZZwqHC1LG79H3xEbd0q+6yWRe0svMjSWPEbaj8uw4LaYOLF84MffX+p2
Deob6JCbzznNrZEHqbheZ6n4w0k+yF5+a+IP9FjYQANOsNxEaHA3bEQrSo043fsa
b/vZAobD9xRFeAymgsTvPpHflw2Yk8964nRTiRUdTrbzGVx2wd79tpoK2V9Qomlz
dKR3NQCrY5gMUiLaAsHXhumDgRsGg4M3kqsrAjyf5UGHUK0MLGGK5rxaqPO6O9Hp
FPdhB/s/FLbUWt38qRpqS12W2JQn7qmJk96z8zn3oBS8KW23v/vB8/UMK2MmD2TV
FGjkuCS7KutX/POuMlh3resgx3/g9VWJi8UXey7nCXdHZMElmqwIPuZTd63ab7Wg
2TkEJcznwfH+SuDiOJFLUcq7hRqum0zPM4GIYCAvqpr5/U1aHSJhWSOkSwx3uUlf
D0xTiBLlNvrlStAzO9gTwQw8LKOe2GCxRuyujgge1+Uo5VmyZchOSuDDgQMcNb3J
ck+Mtrg6MBNU3w3xRRrLO47g8/Gu2lW31sookR2T9YNlbqCva/ZuZrsqVp9jQ8GX
iJXHqH7m6gJCflrfnSyihgFRBeC4gW6VCxtYVHtEzrklAVgJgEYcU7d04ns7ypn+
yesbQE6aa2vjU2iblD5ToUbtVNYdYlNT/k8rAikZlvq6cYdrruxENvrXbpIGQSlB
QXuBKK2P9O3QNcUdFrwIiqBF4VXE5t/dWHHsfqlW+clM+v9NFeAVURShBfvD+EeV
S8DQyb29TVR+KEYYJh6NL1ftn2xDiyCEPg38qxOVhSBD/HJT+E/sCbwb8aLgqVij
d/45any21McMIopfb/KHXvwryBV+5fC78zNuc0LyVef9EX5S7OkJNfyqiZLBqrnA
ZJy+XUdXFFTLaeQqlA0fZ8S2HgsAfFQNYcQE9/K1r80dVfBNvReSjkYbZLS4j3Dr
midvOxWMjuE5VGvdQrerHhYQG6SKOs4pwlJcWeKvbE+sp23ycDKHHZGZz0E8DB7U
SmJikJMtZj7h7e24CbmTvVfudsS8KpFDnNm9ehvL5zKxreItlCMJKtysoOJ7Pm4N
CgZHo3JNPusZT2ld0zXEzgEdobInh2UFoOW4MwYrbp0WoR9WoF/INbI139dJwYbz
u7I9O1z6oaRXM7eWt1iwTAx/kx3vBVCaNNL/i2z1OiKYIGBL7dXg0PP68hXjf8ig
JgFRPfpS+fn26NwSXh+9MJsPsNNz5kp6B+nJGZyJffn0W/ShIMvSmGlvaBayOVMG
nAB6fGndJwgDwTCFFBdXdTVFS2H/l7p7Nidpc2up1gF0RF9DQh7geL1aPBaQ8Zaa
y3zLm1ZBc4xIVCZ/NHgBEK+ahRTGFJZcTgdigF5xvougXQBpvb0YK9d+eolqYxkZ
eQe8DG57z1ut7oofAdJkz8Tzi3rw1+VOJOpeivNBSzhqhGH8EAIlFnf4Bwvq0v8d
JWrQqY/q/i78bjkcDEk5U34kDKN2AL+koNzSygYji1m+oNfhNHlDlbmsR7QOwfvx
F2kd8D+3u0QePNXd8D8V25ep3Ms9RpRUiVuIWrqQD777VG9tJ2KehZGvXQflXa5u
ivbQtJ7M8uHbQoc2mb3zyMDeqb3FWWziT9o7GyhxOChYQR0SCfz/3dfckwmfSlXy
+4BzuemkjrBNKg3+tYmaGWdMhBd/rsQ+CqoSUnUich9Pq6zW5yZwbMMUeiWXmPKF
Wa72YLXGQ1Z30Ya+w1MBkWxr7BHz7MkidZDIU7r7Inob/M2ldyUbriXrD1R3EO6S
03WS4RN/38ibeKCq+rrVt/WEYqnsUcQsDnee0XZ5rDmjfFZEeLNa4GA/Bom/PvWH
84StYxmbCzVmk6iJyLBrgrTy2jFE6rKdIrLYy70Wc6PNQEMZeUXw2rkIfluGa9DZ
zV/NZCiPo6XmSTcEzQSoJvVRcjzSlhcqCpvW1lY3jdpUtFLIwBPK0RkRTyoeTp3Z
nCIpxyRuEHW2hgnJ1rmR6rsvE+ViPCDz6qyZ19gAMDfQX+4vMxpOn+jJk+7iP0kF
p0Ci5n2yqaXXULj9oKNerFhfpG9pA0jX9gNVXtELa+52qPSTc7Y/yXzIUhbRr9d2
gjU41N3KrPz7cygfjBkUraEZKzktneYKBspiVoRNJuEj/Is7dTvOCy7DzxuGzg1R
1ZT8sbKDW3tQMBQWMHi321qKEag7HEJgX2WtyBrbI8EsLsthqc+Ve6gjehak1x7w
IyxKmwSSqyTbzmIsjKp+PCpR8AIsnEu4Fe5G7MIa1tfFH6l3PBjXNBTJILyub2zN
nAl9jfcdNqOl9QG3U58tLNujjCZeXJoNWG11KfuMEfZZVJ2JixV3IUhFJqymkHFq
ufFjRD8aKKjuo9RtMa7SWpxX8Snz+8GXWZDB6iizHAi1yjkQGdMEIAq9LJ22EqNw
ccvbw5Y7YN+vS0IDd0lKwL1XdUQYinE8g1GSr1RmuwB+kBg6GmPmzxORVtwD03is
6g9nXXZdelPF78AReU2qsIEv11NWAP23S1zFebjINv4eRp9DCwbJ36bmRUMLYk+6
DoSCyJo+/rFZlAhtLZ4gh6EVUApNlWjE79/U3m+bQ2uZ7zLT03Tz9G8h67pBl9Xj
eA5sqAqaLxdAKbhOe40lTrvcFremFkQwJMik/U81IWt7AQmm8JSEQ2b+0M4UBkFc
4Q6w2PAO33TxdTPMbwx1314I0xauUFuPv1FUDJWvmHkpPxid4WDrQdmiEPU1rwMS
MR4pcupTKcE1UgUMTv1MEtIFVqChKbcHsAq+4DTCgIFhQcrSagWStmquwExaayPO
qztuEleyzIeEiJ66fL6C+gwD6av2ADHem1GhpLdN4ICAiw+iwIGPcBoGPgZaJNto
VTb5bxqJ8EMd42i7ZNy0H1VpYxVnvQ56LHJZanqd3UZVE4iJvfHrt5oqt/jPGKY2
oCLmKfbtsVdwFc/oqISdP4XdAYStN/T4BWirwPEvzsuF3ujqJNIu09Lpm679EwE4
oX1tQ7Gmgg9zTRQ6hHMUAZMjpKbCFQRWsHWQV9dEX/gBFrtLi8wKaWxiFtueSDlT
k9hofPhW3OdSJciZvmLnrWPuZv3yV2mE++x/RUetPsmqNLjA+riwS26AiXywax9f
uY0ONwLbMCZjabUTANRbKi7I5qH4UugqdWzhwfLaZYZ2e3Pej2JvzcWey/4e6XRG
tzIFinNgRtKfUOVomwjftfekL4EPp5IYDwXfq8njvirkXhR04c7dotz9Z0F/McSS
CLxe854+VfXW6VOnUHFaTisoHuarVDVBvVX6rsXIoPwPxjWhuyPQih+y0Irghs2u
zWoBtusDBcix4+oAMVabnKYPHZoyTgCOQt2DefKusxCUL8kljZNYhFssynQBcqU+
XEhS4VdkCgPJD67y0VIw2GcGIHqlKdI2BuNzONite3o4y1IBKlIWkKvbLJNXE9h4
/hxlGzHbJn02AFZ+uJU9fFLgiIRfsb3KSoctwHVb4NFwmctDj9MvOb00z0XTbQGa
NoeQEMFlQRlqEwZuQTwjwfbJCr8ydmlw4EIezEcv0xqccE9TMl07vLW09BDBahgC
pYjPn7oEIk8UsMzbKcdwupXdYYJVsjNZO4oI8sFCZKc9OaIYfDCFADShrqh9n4ah
QFkENL3X9s0apaq1lYCIGzAOJvsXGF3wKDoCgl6kPgzig2Rb03Bwk/Eu0Vnw/0yJ
ZEQQ6crZX7dNpnqkcurFO85maWTLqXLLrUG2y2O7z3z1/e1X6Gm020XW2FedQuYc
VK35kjowgva4Uw9b9tKp8Uepz9hiclN+VIavF7CGPcC7OAGhnm6Pgtwf4WFB/N3J
+ZFEyisiLxIGX3Z9o8NkMFNQkWT1ifLykID6YYLwNjskhRaAcST8aFnFKKb+imHk
jDr997B1GJxYcwLZERqofMwHX6KHZxW+17p9qXqK6bkqeYMAN6uxPZ86g03HLWXj
4uHm6Etiy6x0k5mjSchX+NO8VlBCRzIMEcXkkzOzzvsRhnwhOur5eIAU7LVfT0/R
zSbMi5842jqBVzZhy2P7UyV6MiN7U1LzOXckl/0c9MOQWKtr2DSAuaeViVZFPA9Z
LpAcRBqZfyZtVcJ5CCMPwHBNLjXBpi0zahiGEljGRPmAFMVtivCLcZRbaTFoT4RU
GTAL1ytml1OSCszvVBJ1q1zOggDVk1BPdWOuKyENRuT/sVzDSkSOPT1O4nYQwqKO
+2jrNURWbCi5yks9SLo1iv4UF9PBKKJiSAQ4kEAbMYWMvQrH1TmzM+savoRi1/V6
Bo+nBtFgJGYfulOjS0RyU6XH/lc8oydqNkNf4tR3LoiIO6NTJKxIpJeNu0OibJUi
NX9c0r0aCsyxdrfPOqggdatQOnIiKbBZSnlyogGFUTFchIIJWFb49hMVRFCW3pI1
UVdXPFcrdzbpN2wWrSr/ssVQcOD/bnwFCobBKzDZqeozJuRQzoovCNwq2KBzgUja
kGjQaLRx78YXC25M8/1F0eEzSiHMMHIsSUXZNMvc5/LyDteBkgZrhoK7qNhBru6t
7qrZlknXKpfpmRfxAd0u39dutSfILULL0TuuR0VEQ1/JTn9mno9hngW8OVmC4Imi
lLYaHMqmlVseL7GelUVCsaypeoKTFqV8Iig6UTQYEbgiBDabOFnLR59O9w6TGnIv
ni9y+FKsePZZ/uMWcTrW35HayVmCpEWWYkHPyaiWXvGP2FEFeIlE6ZZs1FY1m/PU
7gymvNyJYIaGn+xotW2cjby09Q4fLsYuEiinRoBRmj/ClqPyRXJeK1BfgYp05LhW
obFxInIi/lDYHBBR/9VNT93fk3TTzDtzY4WV7Lky4sPPzFby+E8TJNoJmzM52/TO
mGAce+6rv1b1Bby25DD6S6sgkUS0oyv0R9ZGIlL4oAm9i7TqQU1+XY8wjCwLUl8f
d5QYY61+7llOBDiypmGyQIjvXnWg47CNEkrbHrLOiwX4cCYTVrPAYDgRLCEtmoZz
O4MM2czN6pVN1a1w6Rw2fwFYq8vefWOHZ4KuWQWO10ZNiG3lYRQAMjkaH/37d6io
F6rA58ypDCfQExFrUwRDjyo3yYWBziLn7SgxOaHMINhT4zRvPQs+FX8yg+se0h2w
tg7WcBt1aESTv0NrHYEOE4lrH+FgDROrD5CqAzN9y889IjQ06Pqv9HphiWn1h6IT
fgJmPBWhmp7w0qdLmXYT0vITXXYr72hMlm4Bvl13KSaA0qRIJoJ90fcsVCMsNy6P
FrMWKjXavpr4BPTMrqhvVBbV0zmgHMM8kYDHXATKGSKkny3r53FynaqWJ/HYf4+C
/0HWY4iK6ae3ATAzzEEsc9dzPuYv2xoS6pn3u/+BnMZ2eFvXVnVqXPCmVqwEOpNe
mpy8e3uSq9P6HP4iwfpKGSrgY1FjCSgt0Qy5V94IT7/5Doj65Q604ZX95eTBKiAU
i8ByNP4UbqQLxF9D+foik3PXSYFfBYgZUJG5F+bi5/pMHXgyjt1o6Plr6uhli/7M
gijkqm+lrYhqV5RO0PIRFrCTnbe5Yuo+YmJahowWBOrSWL6TlMwF3jYIeI3Jqhac
9dL4h9s5dfuDoMqsDCr9yaeCq8B+uUN0Iwl5oLYZhahQY6SGzBcV5XrmyI+/eiz4
riI9rUxHaSZhnFRnPuEnY2AxU4aPC7v8l5eM9m3mMAQOTIzhgDfBkbSPlBChtPwm
8vpOZJ/irlyd3xjWAxUnTpT8r8HiHAP+5FJ4ngnQYG2u2X01YkNZmkwf4ARdhlm0
/SsUPQZoqXlg3tjw3aR77lvJw3lCsCM5yoq/yMCpViAgofsatzaHy6PV0wO3Om2C
I2hK7ghVgsfRUWZ487YlYDRjwq+YL/4D5LzkPkf+TQ2sdiKZRp5RDipGkfd4zWvd
5frPDLM18mSLjYDXSbP/20cbdTyGp4YGp+UimjR+Pe/RYwQvQ3sXE8aISJZ8MlQu
HKYMuehO0WDEcpSle0xkRjGPJyhxyWIINifwu7QknalsB3Zvatl9omL9v2jwll/P
xuWIuk4r1MIO5BivhMkXi66T77uNSXHIALXT0UkML9MpnjMDLZAinZ/NfnkVXb9d
2/rfHCzhumu38tnrPTYtHsEkuxqGrTRzg+1LkDQq64jalaOw74M962DnDOTpQgPL
xs4dxmepH5tRVEfv45l6YAJKNgzsHlfWWh7tKkjDOMrb26UdTOaWd0u0BSyQ1dwp
NMpWNAuLKP51Vr0Egv/3D+4JccIVOKfMaJgChySXpMAXkZ+810U1WZ2UNU+BHFZT
9bPO8Mk7BGdRCcV8Es60fuW/NjD4OELd0cNCEnUa3BnQqxoIOA6v51+07oUP7WbS
rwPPVgBQ5z6bZB7XfMDb15NxbRpUnO8HxjpwmJnfgfUSb9ltnJPN0+dcAsmdkOQI
5cKJaYB2Q99Srvq5UL5feV0xgdks5ZG9s4cwIMednvG+WjM2rLlxrSXTjE31X+bg
RnqC+MX9C9FgEOiI1Z58z8NZzAZCz7dcN7gXXnu7jYM6GtrfQUnsjm4IdsEJshcw
FhrW+Pbmlp/tbuRcJUsXZOIJN7xo0odl8NwvvJixdcm64AWLQDRx4kWhu0ADXcFW
pfU2gaQzI1hKXlWsj0tlGSyPhq0x3ttavn6RmqEiQ8+/JrL144TzLczoOVdNY/SH
lBNUlRJhhIBMR7Nkqa7iKgJ7H5X7TE90t+rjNUu5xcmvbHabNjVcjtcNf36jDTPl
ftQilkNvJF9ALNItDCpLFl/3WOJD32WmCzf++SIMEYNVzL2YeZuUEubWnQ+zA9tD
Ltw05I/GHsvt+ce2X9bxNEaWUs8LLCPFVoztdZhkW/6Q0VkDc6nM2iZDcCS5o9/B
bU0hFwjsmqltvRsof/bEz+8ExM5QW84c5oLm9wVm2zj8f3PduS4Avg9u90SxWuuj
TNGbVHm5vZ0lCMPbV7KOO1HptWgjC0EtxsRoTpd+xXYC25ioT29vFCFez61QnMIV
055BLwwAmaqHgoHW06khHaXE4GPpcZTXIXGsgPhM/tS3o3w0kPYVy5FayT2q4RBJ
zDqtm3b1Du7agOwia2r09YCW5oXpRPi/BG3uhjs/NEmM6lzgVPO0vgYXkaeh7bIE
wV479DTzF8y4FRvDiZwPKKq7HpjN/knEXUJVnlzrchkedsbA3InYYYBnFquwe0l9
Zd+9Lpw/3K7gWzLjPpHwYe2YlJsEsx+cuD13I6Xm1Yb0IDWnTIDSDHRlp/ZtVGvy
8mXlFvqxqlPgS0cuVwA3GoftVDqO9e4fkggDKxOFn3ZdPP0Wj80jJCiOTQ7cun2z
Fo1hS2JVmbRJOGiUuLLc4hFQmX11GraGdy5k6gaHzFDd776Q1JheNs2uAIXpJssa
E1RU8YhcolVWB//7VbbcFxc74c1B1xYIXZDs518r3EYxjndWvyy/9C0zWtt2Lm1X
/YkZEcHBLYSuISRwy0l/i0KX3lBOoq5mcVlRRF9iC5dslpD7ymbprqB2exJlNL/I
sXtQWbLGqoB66vlBCdhHKg3sEjLb7Wfmd7Gx0Um3fWdDGp+V2WMttMWg6D/rKMp8
1B2SaU2n38quqckkA4c9ywG4RvNtNKS63kDeezrdVg8BE+pgL2HXI8uzZjrXH3kk
COS3Nzsd0AVY1j9iqXrC8+z00WY6PwmLOe6OQEaz7giV7wu+G1lVDPNjgy+mmsUJ
nZ8NppFKvwmqIcXpNNf5hmMI+zsrsLUqNPdqYdHHNgYiQ3lz9jtaBo7DSSefEN5h
9NZa1tZe3hwwzktFdg3ameQtTIyUtRdivCJOzvEkqdz65lsbh/Bo2h3OdYxipt2e
j7Fid0VRHpOvDqnFY4vO/QZj8sKZxury1jK5lLVBvEYsOwWsqxv1poJCwq3sHIzL
TjJ+Er6Iv0O8x4bQS0MJPwImx6ZluuzWdzXM8xrnFnWTTyK7ZVx06imwNaXAzK2u
f4MDRMLeMJCHg5aroQEnS7KfSbAILJc0QRwvTv/Zt0s5P5eCzKvhrKKQOrMzxzjF
duVxFSF28FuosVtlMOnmSP/7nZ8N0HJ18ixauRUKKe6z6LO1D3eEqCxnmVxK4ehY
DLZEpWrukRWQwjg7uLXak8ZtholPW+MAjdxiHctdoAHUh8UzYxC3uniGK5yDJjwo
vxlWOZ/gU07T/AiNwQq5nmGpoqFBIh6owxLp+Y9rtcrHdxf+BWExJfsUMQr63brg
xtrXYMoqqr+ucQuVVmc2z6rfUMWNpFU5d3W2rFgp4QRoxdhR3Aq1WorYcSiglz9g
C3Xye7+Qh9AbmwDhkUjSWxPzJxxeOhXfIRnCe0PZYUiL1fa/g8d3QHQmUmaaZyOZ
VE85+u5xxTKSsD3zzSB95lCIK/5PxVQYTqMWBNKcS2zTI2kTBcrv6i9nY8ZgjcEL
kdeCuQfyCGxmGaeWGQ3ZwWGekgA83k9OdYl8D4Doc+/NVpgg2MrMxUP2FiL0YzJz
XcGPIcGJ3ewdfSjWZqTiqPl9VqhkGgmkQGKm/I49xizau7MG4xz54KptldC7bkqO
8vJZsDZc+n5rQy/dNfSx0f6Tr75wBwfIDRHhy0YmsvOpSopucycEcnc8Bo+REHO/
iVJqPZ2QobQe6En9tqmH5uXrXBTHUc8dp4DIMYpgwZOgf4ulPbTJo9EaZHz+L1uS
jRCqEW0LLAJWWZnQJjbmFvj8XO6RUF71kBDGmwIc2+Fy+l3FAcNy5LGVeD7Kt8uc
L8/79W9nPoqMRFHGvyVUs60qLK2BumZlZzhj3Eynrv8zaGOy9UxtFxNGfveYxlkc
31M6YTeHGz1bdhR8lNDhFnwUuBwoKICtz0NJBB7lxKzSM4h5R5o41RBUdoIuJsml
vsUkLgtgN9YYO1n2u+dY8KGbB761aqiwoGUyFWLz9ghpnckGjHueSa2kH8rT9wJs
eJO6oayIWqosyRDSEoYnbu5SJ0uKeWN3lrll0tcLzt5Fg3QvBE/rpUrp2AWGJZEI
tlg5LMHjeNNPPLLQJ/fnxSJBjLOssEy0YZ/+s7tLc9InHnwNH1PqZ76k1m7+GYlJ
Xukj2mZDkLi1aWDDTPXRx64zNHpyIhr6At8sifWajDzhTkxuQfEIyUBXZCGVgRU4
61FWFyBvF8bypTYwxj2YkDwUhqdco98LeaXjOXhCZCuPq+WzpEUGkRdQoUNBM/zB
oC+Ub9oQyM1V9Yao3q2EFupGzslq9NZj7OG0V+CZ/g0b+8l+iyvFeupt+N8Pf02/
sfXKqpCg+kubRk440C74oMTzHGpIdwh6UV3iLjZusGlOLeMTA3Zh5rkc00c+qAN2
tt+1hv+Zn6q8Yhge31SMmccwcGQsVaAPHhN+HMptp7mUOJWMQzF0jqGO2EAkroxx
JEMIeI23qkwlWnukVqAl8EgBP6pJX1+DJSO/7T7dvm3BLe9nYYYu5dCpr4Zq7TFm
4PTerqlEb+nMXHgGV3WMgt/tIUultEwieNmgUTTqyZmL0/XB+p9+PSLBJujTfgNK
0YmL8xjR8B4ekzzV/ylQ3pVHQuXfRA0EuWzUJk+BUHhr/nXYXDUv2FQnDaYMXLjO
Q+/7YRnZX7LXHtn5Zld7bGeiXvF2HxyiqkpLmMXctVu3t34JOxhX42Z6csz3F9rl
UiNl3uEkAFkD9Vx83XKP1T3DDY8S/LkU6PUD7W+3FkFzo89bKa1aDA4ZB2kZSQFN
IFtZmBYE/RrWWDSZMa+yU+V3QfjPEYgB2NWxdSDI0CuV33/dwlSmnsgTArO0YTEV
qyPQCEpiAb7WPGoIGevwiMX7ZkMYXV+hQrga6/TxacWX70T+eo8t8r0GOVwlkBA8
d94wZHK0TbU8irsxMZTw0dBWKHURHfZ1Z1jJtvyUnMztHH7vdcW+PxcxDCCurf0r
xucWRBxMvvZC2wdhqXRRZ8ilWiB6Jr3ByxImHOY58n3qrrDbMpUXCrKjidEno1qY
h5eX/rwmXZ+3jj6uJY+5Y929H16qMpKnzdudja5g9S9c4s5092R1TnVz0Ra03jz2
TZ23dU2KciTOhLJ0TK9RQPK1g4hJNFZUjqOn7UBtd31LyMMN9nvLWr9XaC3QJCHd
2UQHaqsde2keDIjWzcKmY0BXa9WJthXmqKD04OKoqjbAhI4Zu0Ke/if4av0jWINc
VoH/M2tyoSMeufntybACyR0zBK77m82UsZlCb8+RYEp2C27nK+oB0emJLsFo5qb3
AicG47v2VHX8SoPxIPTHWhxFz8JE3qUvul2NNCiFa/+KoyOoShJeAUfkSt1rY+1I
kfrHn13mlEDEAp/uPPJAr1mApf4r9dh7+8FR2gA1OsIunpXW5HiNI0zmPd8Fcn3d
udn4fGdAz/s6i1IvFBMwJxpcooCFBsBtLjTKqbG99H46JykIokc3RJV4UTWtOoaS
+XFog82tJUWTYTBV5T7hLcWzeETVF3VDEKj2fZ10W5qu4wekcRU6Fm1rVGe/t8UL
+pixod9TrBan8HVqFMc7j1Xv+VhJz8dD37fPGUHqIKMsNDiHxqW0gfnQzy+6uf3Z
6bbxCpPkq9cOQW00vjFXgFuyCrrt6qAux5fI5uEszRnH04XLNHfMly8NiX3GNGUO
bu7B+rParHJNBjVYE8hRVxs05v9+ANc5SDcegfmgkxImUujXbPkZslI0lia6jc/z
xgXct1Nhl+GGx5aSelbHvK/FyXua8rABu0M+CKNqe4/3jcfIeNXRcWhLXtj0NeXQ
xRPbrt4O9nEnKC+NOzw0gcRqpYYx7EZiZ6r7A1C9Y3vzlFfj9Cifnfxo76lmjgsQ
Zj84BJ3KWtheNn8dVuVMbmp2wPHRpi1vr4V4ak+kMkO1loPixQD2yDh6o3WLYCh5
fkbz5LSTdqBFgxRo7EPtI83dF9pPLRXp9Q3vmSodZUqDGLGLDM3OWdt+Jtirvp0g
Gfv82gccQvOXtxjtJHacoodWzBCy46F95Z+de6x8uMF/qv4W6PWufCjspN1x+czj
tiWpgSfVllKyInREVGYVHSaf2rSxHHCy34Uq9nG1BDgSpWE2R1fvjgI+inaGAPM1
OBMsMpoqJQZ1AJUjdZoO8Ww7GXc8TMVjpfIvTW4IaTB9hg1VB3HJF+VWCISsNss0
Talsb/m2f8crsKquFnPTqJLR9mR/Ja542OqSsePpLo8T0bs9YBIPJCK5WNAGEqUL
hK2l6leYiiPPYyTg9rUM0yjKrKXCfWywgTDNSj55UijODb3FeV0SomaWWO7tUF0p
96sxeqjFXF/+R2sBOrbpK0Pv7CxepIauC6zJC7R9IfGtgVqMfyEQK/jx6w1NKS5w
oYW7RLLIXNhyMqB+VS1LDpQ9O3JsAT4MkdVRzHy/pbAvVjavAPM0Z7iBHDYELTUI
ExMrdK9OMtf97XN/NPUnkYVGorVusA2x8eD+Rbevf9QoQ85eSyfXQcjCDN5HOiIM
7oP3Dh3HB+PO+eQGr1YSXCe/JzyYcfIGshQ7hBqpc4OAjwO5Fwiu2iEagkTaYlxB
EEgSPNRM+fQxqrD/cPCmL9pSLsda5p6yODDQVIMFy7joGaBOwvQ1h3VNhAVgbahr
ODJeu8b9mTr7rJF1nySmm8QrQ24r+/uNf4Ez24dW9FahY3EHUboY8ajvdM4HRJRu
BS5XlDFcBDTkWw4H2hZb9KILAxd/AFj2aj7lo7BGEbgSm9E/iCoVEtehsj7NVdSF
PiO/c3jH9w4GkB6xFTs5PK15jxaN3hTQN3DmtVizWuPDagwD5u/xG9C1S1bdRQsz
wO4WAVX34C19YJyUIUpudyW74wjD2QFxrM4IhbgzCgQAaWT+phuYa5bCbNrWyh9U
rYygPAgLL8WrNJzkyILdT9M+8YC/Bje7JSWEZcqC0sr89FH0aQ8obAmz56aPLpDn
egvTAHr9U8bPYqawJglQvrJ+ffhV8/n1/zONVq/nq7PFJ5AMq5KasUx9l99FK2AM
Qv8E2ouInwU5WhYnCsBkxydtvNFkCKU0zOscrGCuzMYjkI90MwpCCbWHcrccA/20
3HPgtcw+VpF9fjgW7Hf+MyNAFDXw3wZ3oCLPN3u8vxMycrUQudU6s+PADxzqBDEl
CcTdemvzbpuZ9xnFxUsEf5clSMgXJSw1+M0/4cQWUbIvfjQKHBzc/CMEcV595U1/
hmMXXtVZT6k+Ye3anImxr6zHzUMOQgb2EN4TH5dPVanOPeoVftjHlit3oWJdPZsu
7nSsyuPxcmWfwho9FjHLTITbbnrN5NPiLWH2ByWATxrcC3FJy67mEPAz5krNMZzH
amqtovA+ghpVd52diUtnAkz06N9GzKzGIl8NMN5WbK0XIab8cO96UNGWh5ut9q3A
rdF19cJEV+NhXLOcK05MkW2ufBWQjmP9oqjzfhXtn83NTgKbSMOaiWeMwePy9RDU
j4JR/4y4LIwF5v6BDzVYsQnPEDG5h0OOFC5r4YJEYOdkSBNEY+bUNF8CXxY9N/6Q
UbWbfYlikj5QfZSP0a81jb8rxM66wnHN7y6pVHmDG1R3tO0dZ6P+5nMo+ItxeFJn
NM03prFMyt2/5cz76OOEUvzvjzwUQLfKalFHXNT6EaJrmO7PmD76vuF8rgZAEv4W
MEv4AdrB8UmdWPnQ+/YMyakFYwnBEpYuwJER6t2dPW2kHCMcHY1R38rcd7kEpQDd
Y/lLdmlwubntCiuNCbnNPg+dsHlWI9bD3ywItW9K/1c+CysY1S5OOXkjcz96wbnS
oKr1u5jjYxisPu+N+wulbE22/aZnuGquMvyxperjiQut2wrZZoJGad2f3KxddrzX
cOqHuI0+fKvPAcmOmIFRWavVwWyFurdW2Knl3u/TCO3qEmBULcTbVyTO0GnSqLiZ
EsTBieDPBUkadMtfVn5pemQ3LSRk/x2U7204waqVtnvV35+E45i5vaHFLF2V5uuS
qZLgUThCOI5pjCH+z97QmAmQa2TET9Y+CsZ4BAx12DpcRMZ1WlOzCWgciIEUWP8G
O49I9rsraRo3pzkoaPaBrk4aRVbhHyksshQInKl3KyJoaWYX6yA2qTh0SrdHsHWX
oBAeV0nTYuvDZHmF/AYS2+qfri08QiR1H/s51sdxOzTyAYvb907ladMqJIll/Psl
7ySreFeTycJjz2DwEgefILCJJKo2nW2alLBvIaBysPYkteqwyArciD6Pc6BB8JTW
ZVy2IN0RNdgnqS6S6agSRpMkfBc9LhZwlUADuLMoV0fIid1cSZLDlot94TYe5G6j
U7y58RF/rc/QunYVwjsC8g+HfCR1SoKrhsnTG0QPGOYFy8G2MnpTW/lFODUngvp+
7cihimOjsHBPiCut/QiM34exNf8bJhwRDOZnPpwvdaXBclpakfw6Ws17ARxw5LaC
6Ofa4QO7rQTZU267Usf+jLbAbvSw7ioI2xmCUhSaSkzX8cHOq6GGvkO6/bxT+qeZ
QhYrD4i/THXLSYhnKQq0eQh8csDKAbzR31sH0qjlbYVVsy0THcP+Nv4cp2FI6CsR
ZpC++UqZ/OtEsXjNvcNZ1ur+4GE/SUt2MJsHs6haPE7LEPfXFKRObp1Zqcneeu7y
Np4P3V+8iZfmtp96ap3oFSVoYnFu0ACq4WkGN1d3W2J5wvDOZqz8fOCEq4eX6pnQ
fCEUGLSwHTxgV6arj5hRgiriwnZA1HNj1J4MiXh9CLgmnmAHJK0aMki1EpM3I81B
5mIVfl+hBpC3+GRpP0WmScSA2bSQEc64f0aycpen/U3yhTfwt3iny1Sn0s3dV2PQ
3LlOghzc9NuhqVKYopqS5lu4PbdUO/U7kySIgyxqTzW1a635oJbZmpOBhulrMiCY
7eux35ROhXes8dmV+yx2F66wzQZC9Xn8hxisISibVhyyrNsjEIUpdJT3tK98WQHM
fiJvsmcoDsSjrspwxwH5+b7kZnGCv6BMH/6gszgAA2SWu7h948nE+d4dMqwDlqYx
Q/4FUm5ZOCirPWLTjVShOdRKqzkKaz/srMoV+t6lcYVuBFmIIGaSzcepeCkYcxm0
1XoDLLO5LtTds7UZpA6oRodfSkHQnqAG/XaLnP+JIMTW6gmqgr0VUkHU2tEdLWsm
vM/4tS+vfb1twiRBenvWkBxRR5KNv7jCwXqqGsBfrs0H858eYZNSwx4tFLAcltNU
zKXDdLrKKC9xMyXZueb4PfXlTd39ypRQXk0FN6mjnamuVPcMyI92dc0evpv7xl3L
79DiihU1ioSm5iuFm5O3V5JFHY5mlIMCiX1ncVQWisHhKQPVbcXosfcGytjzulzz
nW/oljUxLN1s0mxr569G8iBut3g1qUQROI3UNSsoSnPzEFyLrTuVBrdoXP2SWw8b
XUvMyaL2RwuwDF5NH2ee8OYOdD5oBALwO9fpvTgy62AKHyUH4FYea3Vei+WW8s0J
vu2lK10B7u9rIO5rGxjqErDLmUMBJAMULWMYRzCtRBrDzV29q61hQn/3ZGwEE1wB
7Oj9GpfdaoqCyhKpGQm973G4V0haWjNCQqsbo3cUCIG8n3KVkRrTRtibRkNVFBq4
sMkfyuroyZQlprTfBz9GKFrUQ3qR0bh43YKQnZUlfGwp0QuJWi90Ka2hWXxGSCFX
9xRNfkALIUofERczXfjpewgCRFL9Vwe+eWzp7JreVS7SN6ZTILrGPRaOH9hHYPt1
z9HRhPyMonxmY71bfWxbWEsUnwQBbpxivAXltBGUb9aD3D2dACRrx9VTPhwMWQFh
QYVYoEN8umOzeczVNYqYmUT5j7AmpximBwwGI5yATGz1ygteIfxosUnj5i0rIPzX
ORJm+Po7GERn1rVdMc0DKyJP2qkPrN5a8dlrGsVxs/SdbTSgxCLihIMNwG1WqzjK
2JnD+y6YHM5M6/0Fe9J/3ykK3rOyeBM8z9l/A0VdfC22BSpgLS0oaf+JW1qKvDck
6bJ0WTUGfmuNNBW7K1NNX6EvKCTtby+MPhjP8X3YNyJL/5vB+ROh/8UTkRYFBN7s
/SwVHO5kC9y7+9R+tP8Fa2rjXkFGuBO0/ReY5JpufSRcACxeKQLntL+EAybf2x0p
sNmKrUFcaEv6oV25whf5TzH77RpoBMVAr9mYyRRT2ozJgOSvQ19uwCqD9U3kjPsS
9wKpGlzUy5lYit8OjkFWqgOCo82HYUVikxH9Yh7HlO2f41P0PsfAmpUhDfc/mvn0
OU5F1aufxNSZ9tQj2tgfIrSogitTELoyBNn4ErpDZNgm8MsDieULm3EcVwnLB9EX
GQvxF3N5MaNDAHbKeDZkbhJ9hyOwWI6LUK1ShFLTPckMV0DtSQGyzB+kyflhQx99
badH+cpLRxT1Mp8eWqq9OoWtXTdIKE9PeV5cbByHUVSlfAXrQfdb6N8H50sR5VQ+
lWRghaLWqVC2gx/Ci+UhIYQNiOCjAwwnxJLPNi1OgORz4edyGdau+4qbOzU/P87d
njKQV2gCglAoOkwdk7cionQPyBPN57RUJhHt7/2+suqRDl+LO8HsF0hcQDhzKcXg
WX3iaZjLwW/aotjtrVIvqyLbvgjHy1vxW/quxZzS+3N8SiephmvQ5j9dfCtIxTNd
AnmmhDg/gH9fLthKfqMgRUYUXGasJw+ooISHH12M9o2vC059xT/yN8xtuL3XHd6S
XAytlNf2pf5/50r6VjBYUiBnA/0F5OYtqCwLLyJyi5OZWt0XkulxpFFsS7l/ZKtQ
YRGc6T5oVMNEZgrPz9OGlbNTBE43WBQqaIZtrtXSb2KCj9lKSXlsJbzMMzqlMZA2
MpYMqic7tH46aq33RYgFuYDm8WZXiy9SOrZ/AGG87DECeZv0xS+usgj1iIuW3DAZ
VkQhRxdwY9cLS72ZJqEEIg8HHQjwQf1wUmKS0frCwrhO31o0jTW5F8A3I28uIimg
Yt9b6IEcWg05ethDWTHa9wuYFELjEKoKe1Lj0ebk6zBMvOaQaTZDv4HZpb9DlDMY
+6dlCIb/8G0ED9OsI4I+8gwSY+AT/IkMRwfujn4OfAre3lGtyONNxqsQSPUbYmol
Z+pzeOPy+TW/6AJlnkV5m4rst8Zv4wwDNmudW/LWttiMRhn6wzh3iHkjsSTonuBj
KfSChP19yPw3CVPCnp+OP3ET5Ihy6QAoLyzqXVyGHYYHPZ30d8bsqqfjXRCyfSPN
ohh4xY7bQzn+ht/rpM8G5gnVy8gt7J0P7wVqOwKOAiBKWgeHO0fb0g4IrJ2WbjP2
CP/YAsMgtDe2dGVeGPXdqXHXFDya5e5AS6+q2oAjUGgPy+Lliz3SWHqKFvzeiluE
quFkPYnMYcLQkw4kaXG/tZGGRDGFLO6D7lAcKrk26RwEAwDfab4HLGZalBrGnNSn
7mlx3wOSFHBS24unRZAexTSGD210WOV2eIktSDXX1ryn0zF4Sv78TVLCeDgcwQcm
MUFIYpBsKKlUOaiEKtG7pLsrY2xGLK3PYRxownZV5rcB622ml7afHbK9eteLoRu7
BMqB681hIhpOy1CUGo9DuKXbRIgEnZrwi72JK696tsTlqVpBaRAy5hER8m7jglLG
vaT200x0Mlp4UXUUuuXXdWTjCK7mYjgWOZyjlUvLi1XeGSK1Ko/cpn5N66Ucu4Dq
8CjGttk7+zvwd0ek3f+SPdoNFkrZ3cC02/r5nPi4LTmgprtom3PBAnXUHT7QWJE5
DreJ9KW+XH5NcBmWGtzI6GniLmFyNikuWPjvRLfyAB+6PhYKlCLp6OhXYV88ipuD
F/bwItRbjgfLzsuwna0SaRla24fDokLLyFLGCUFJYUYaqLoCrWmmDueqFNOiXdcj
uG4sozpNI5ENju7gE44/qF3cWtzzfug9wroPjCjMygJvS6998i9jLfwmc9AVVCjC
YatN5RHuyNWdaaxxTtS9VXqxhZwy7N+WCSivLiZLwwtNfiBzWpEA/rGZ95PgUIMd
nJT2ntKfVhZunDe42cVnQYuZvtwXEhqhC9fAQ7yPa47gOuxsKj2nXcYb/C54RYJ3
sw43qC2VCwQVbe14ANqrmCG/8esqSNmBRnx+cJsH2FoTW9evJ45it7ZLvCqDx2oB
LIBn5Fsd7aD2xPXhyDPyiQ3oSK0qLqnyAVLBr1b3SlFQ922mMUkdQxjz+4xuFsG7
al5wG/X3XN+T8pIR7zN1fycHBD2cVsG29mwhIK9YQNsSpe+VNH62EVnP4WI5Ni0f
YicY2nfv28IL8T+eGHSh50kf4gTCugKcUxBLdVxIlMS4Np2j5iLaaWH2VjdH3XKw
HKmoFFPMKsKLZKCfE8HayRdtrHDCxPqyf3pMvsXKqSYpYJFmXQ7rgbzSVtoCprUX
kB+5BVawsXVExPLynfV/PzbiUp6HPUKwGJxtt6veTBCwobtNqjGeTNsqrRXjdOfs
MVs+nKX2uMsRHCTzwckEHCHy9lu11uTKlldFubYyZKtqigADPrLeiY8mXux8LhyZ
4wbpnP8wLhFKuPi8GkOeIRi4un+toMyrJXiOfenyQa1UQ2Z6CB8Noz/baS7ZvIpi
MqvVyuE2it60lvOaKtq2ZzmXtvrJldzky1gWKrzpDgbElfvrm+R0hy8bidOlrFX6
SDY1GfScMbG8SH6wCDhdN2m9ZohWeWE73mFolYEC0tUzyqtlA5cc2AIAwlKaSD9e
1VauduN/e8RK4EQHxcUyRPUQdSqRpeCvDbfBYuTVBW4GIG4KnzwcOkPKgS7BB3iN
0IZz2fcJKGtT6/nckZ5BAHIH3RC1jES55M3JUpSXuzR/IKmgWkEs4/llQGf/9r7M
WJVqMR33QeHJTXV9uXNhpm2Uv7S91Qd2v7prA5UwnaYQffY+VIxEpVR7y4g3AZQ4
YgUlSpkxcXTb4DF7cDuKt4Hjt8Vi9A96DlNd4da74PHSJpM+COkEHR2i9AqPGj/U
AsK3wNZOg6w/Y3vyHlSznZurgxSKKVsBwQsQBgfGIB1G7imXtBHCrwXbMoIHjWWp
mbwEWnbzW+SowQTmqdoPqX4vmOoLiWUls0tO+BFRbS+1B25aunV8eyQ/PXP98HB5
uziGcdU+w8Pg3ipTYXF89L+IwnTPpY4KJHw7F5ti590vhgy6QkP50yJ8XMzYrpj7
pBARYQk/y7t3J1zS/96ORAE3ZH0qIRW11xrvpB0VhjyPoNwiU5WQ3/QTHpLruIbL
0BBcQ5WFYMlRw5VkiZp5NhaUHUaWWgz8jV9O6CQ2WhVnMjEMcBWSMc5spDduypPh
ZmVuiSbLuFEIyKtVPh+khiOfS0QPTpsxDINXVtJBaRciXTdHttKB1JIqqRnuOjeD
QGTnW/mfDsBH2bwl4MVGJ8KNqzJECe+xjy23eO5YY8L3qJUPlCNS4KPdaj7vpizk
TqoBsmrIlUQXyoCvlmO+DblBZ7QJyFweagYcWm2DlqPXKBWE0yGYJ2tJWM4z4JaT
ghTjWNrG8vmw2iWr/seymujZezfyho2cgVmxzwLSt6hjhs1U2mdDIfmX858Tld85
a8CE/IevapeWlZEJiDtdetcwHqwI5NDidJ72M0QcHtmYlVJESaWJSwtTUt/ixpYl
UCAA2ZG4ZpH7uvcOv72blbtWzcUEEpqO/W2Vq9XjeehnhzDGTucsDtZYKf4jwCG5
HdabSEtFsUt87AW+e4HZXKaJ2UFfBPu31L8iWjq78vvbezo9LUMCZ9+N6c8NjyiT
u+ip+QEvPeaJ787i8FyiPf9abAgxotITGcxGTN4gHxefYPl7qR5kktMSayGdx+YH
KGG4FxDL+5M8rELksdBUKjx2L2/H0RjoGrWCdUB16fd19tLIE7uL09cUSWedJHO6
ruknL249G/Imex7TX7k5snO1iSH+rYj4LW28cICe6fpzpHHnXQPlJEx8Huqxa+Ml
eJcFba3pGb7SlwBN0xo7NOX7HzjsCrJ33vO/+3nRXaDxVrmLjNT3uPhS0N548tpu
wGLgFFVKChlogb4w4LgNk4+34eW0b6n+ZtXH2Pa3kvRPOD1BERf4lH2a+ynEpnyx
0ndy/QjlIX6DZbf3XpnKtB/WgYdW6xtr0X91650dqMk4oULdqbYmesX3Fy45/gYS
k/twmSbYYAh68eEHWHdD/nXYyZmWidF7ahUEO4WXyxDSXDP0DRq72h2k3gusHo/O
VHeN0i5sBu060hBXWYN6WpOkc8/4yvG6nvDp8I5qdmZJ8yqel+Whdb2S5fy89RzQ
bUNRs/wjz3oVkmIWjNzSnyoz84qHaoyTALjJWqRfdPczjRyqkQoLaQPzccSRhsiw
qs3Y5elPvbfYEOaXrRrMS1nibWNTnyNdemlS0oN+Pm2nCnOPbzyWTcXz4RX5AzF3
kfHZl2tl34kY2PRDsDUNbSiRY96gK17MMm8p9hVYp+N3KfYglNg3ULj7X91Wn7y+
KjOzuFzYbk5WXzp/eXJtb6hhzjjpyGavHBGiSgB6H11qQ/RFPx8Z08H0qtoYlMUv
CpgZatY2nhyXI/xqzOtkucfIH7ue8e107JIgKFMi5KUsEi71WaTCd9zaZ5+ctzTJ
jny0TltMwM1VMXXIB2xbzZDZZfsRGQLYZHUZ9hoElMOYnQDxNwz9cXFGvxKizbLd
NlwF6zjJfUYqnJlILDQCSG0GiIchI6ht0OQUcDN1aTrFr7RvFDgDfc1DTqke9BPp
xRWe3rgu7q6grqKCyTHW5qqDyVvR+oFXg/AzQaSnlLeWG252q3DZrZiJ46xNduoS
ukZjdjLip78df9t7pN1w13bputx4O6IBZcCEYj61JFbrSGBCq6TUzBQdJEBxAv9R
lTE5MEFJKz0jIdGwD9RUKdRBT80BdXgaqI21/fptluGKbP2+kVZWjp0v5Ler1+tR
AaqY+/geOX59m6ikvXxMp6HM+IhNRbbhLpEhvnFuUJk4A+FhSGkkTYaI5C84Ua2T
niE6OA/vFrHaV8HKHdol50SvLYeMwWc+SHlWJNamHSL7DWS/UFnfwDf8tMnNTK4i
uS4xTMaxnxFotd3VC4V9BSQ6S1tpNPTJXyW96Z0cobMOJR6k3nOMIzTZj4PZI5fW
cMGlYY395ixDqf5Dwdii9U8Zo6HH4DsF8wcgr0mkugrKUW7s45zyPp/sgpRzGylx
OFRWvBN3bbebpPxnR5CeiAiaAHxSFgcmvBCc2XcS/5IvuJhV9ky60B7ARU2gfLCF
dvK+MEkP+j/Munr2wy9A4XMkeV5jd51p4smwhQLRLKiGqD6eIMjRIWSMxm2fpzhy
R4EpAGFhIStARred9P8E0K+ut+jPu1IopY/wrF9sldWSUb1JOkUoBEf2zNLCNZ7H
zmWixp1DJdMxdblvlN4skXwnPtj3/B6vtU3TpxeM4G3kEpVcSGzSIxFUBSVBpLrK
aGLDqftqD5M/2ROjWSGGn/LdIE3mwxQHAT69DoPRJojHKp5OeARJ4rKYZUAlY4aN
RvCJQFHaIL80qs9+ASljUsFEQBtsPNfqcQsYOygkzBVc+6DQcxpBx1r3z1q0Fwsg
tv/JBci8rbwcYWnWfgCc/ZE0aIXhd5rcn9DOykAluJ9I9PjvbrbxINoz1hxY8hK1
MgXA3Jztp695HVKdKk6ZPM7oztZRROLMgBgJKbhkS0Z2yNXvgk58qhGmoMW1hsQu
9ZXRbV3DFN900M2U9sqPIFhAbobU82kQKflC6DsJmCGX2zutiv1/4s9m8hLWJYSE
V/XFIvyxZtxikRn44kwa3LuYS77uqGWgQLnRVm9nPolXXbawigeXK4Ow5Xqd5n1v
XngBWkA5/06UmbXcy7e/jd/KhO8iXTdXv6LBvlN1eywY5T4hvY7jCuvO4EMs051n
CQYQACsiRRtFq/00QZHRfiLtmWXb/wSPMz7dfFL30YYJOo1NADDtmdd9ewNUjs59
yjAk4eh9YV7mC/DvARrAwVQcgw0cg5v78xlXKMSWUe01P7u0XxecX7rnBXIr6Fu9
CmbcPw4G1+K2lRCTnNDNcRB3STo2O9/8av7mTTVzgRKcOsgIpAF4psyzsePnJtXj
H5L7dlI9LbZXjUpgn/VrayFL1AqQIPpboK6A0vMMvy73x5HkhkWVywg+sdh4S4mq
MdrOSaLUlTs/xEEGDWvFu4cPv7g23ZS7nc0j9+eS5KekTEI7bDVmiBYs/S82Fsk5
KPtrrYxArG7L6xUO9lhUdOcaFlu5rSbhSSiaV+q/G0hkJpGarKW8XjZ0zvRQScSp
jLhfDg/kPR2SPPF0qg6XLtMSou+bupk/D7eh3Q3bVHbyv2LpzK2ZHQ+HeNy0GdqR
DwuUviN2NvNhoregDcZaRoBDOGlXkpjmcdbs+zXQjvmgH41vioqyDDy3eVumoORb
wvybiVp8ATLcPkRDB9eVpy7Xq68SC+2oGJF9Ot/vhVaclvJTolfisTVLLkiTCjk1
T7JwiD8N4f2aXybU+JB/lknde0s9tc9srITLMPHPuJLEtLG6vW57DQfiP2tr9eXO
nwMWb+qCHbOrdqr2628j2I7RaXOuKPWaD/No9XEywznfq2dGROwQPduSmikP+Ek/
4OIAw/CGHG+vEF0MsBkE782TcFmfalqKv46hJrX/dbix7f4xouXXoLkUMQ8eXJ3e
+oAFE+Xu0Lqee/MTMKlihjReTk8mb1W0Px/UOTSZyRA0HWFRArNZ8YJhJMAYMNCf
M1hrp0s+e+5jhJzglgU3iJEDBNBWNYfbmZOvqZXB+uj+xnk+2e0tTWqPHjccym2c
mDmm/DUR2/+Izwky1T6gt1Tw4HUlLPARmizohQvsrLJIivuBDwT2dEd1/yviWmYO
fKsZ6RXAagBGSk2DKWGXBA2LIumoBZUVSHLZQQunEms51WrpU+3+g/21CoFTyMXW
iF/d3ypR/nsWWePX7ICDyLi7GeZfMvPaFXhmYM0dLBkeaGJa664vNxL5FXIhg0HK
4nIipexAz5Nmtkm3xl2E1PmTJnR8AP5Lv2A6TYcNEhJu5yVZo9iSZm8hpbE+IGur
DZ9GKbkjlTOYO++rx5c8k/qEGStXTMi1UOY5cPReOTB0SPYjmWqaCK4a2GVZZK4k
cPHvZCUwonYtA0x09qYt5eB7PyEBPZf5a68s8hfIn7kMQATDMkoXvewOzx5h+Gay
VZgh9ht+de2kDPIyTbSSWi4Lbju1md6a81OyErQSf8YyDUiBHOVKLdUSqarzY49f
m1tN0wh1Ia7hskMtFjG17M91juSQBNLkqlgQQ11EvxSmb7C2vOGSCABQCstoks8I
L+Bsx0SzGhQ5R3J9mvkuNVqFIsIHQLa6eaLZ00Fo93gMSBHwIgaKAVIo6WL8D+DG
LbbHblJQkZQLPXQIrdzRVkszWHgH/bkiRQj0WacUqFAxcQ1yoN1yLEVJskhscwgU
AbC40eaX6c7avbPr+jWcPV7LPjZHPQhFRcolPQ9iWgOAmGlWLuGQe5WxhDQ87NT6
9wKHhOgr1Kwbv4uwS8abC+PIzG8YbZVon0eQRakToZQb4eRpCjklELeZm+qsmYAl
tcM4TcrG3FBjiY8PIGC/8t22p26uNrFHTbgtJ7emVofn2zhq/T1Yg8GyRTbb2xlD
M5INw806VrBzOqcRRE1EYqVlhNjKEOF18rbYfQt9Dmz06nZs7dJgfl//xRpaPNyw
zl4CaPuOaYL+o/qimbFwZTNKbD6q3sb/GfNK6W78YLfGYaTgtC93Qf+WRr8P/Rlu
2RDsXnpAfpEXp4pJvVQWXo2h/oDNbuXl/Fnq1J8JvJQhJ0xXyXVIZn/9UzDn2JaZ
j0CYz+lWi06wpViFUXR05EGCFT3ob5n/kiBSSWNNNWkPVDvhxyBOkhjR8/BfmXMN
zSGpFnkKUQ116rNN1dzcr2GjrD7WECAPV8H+2UpAfPu8vMT9SFMWuFSow5T0emOF
ld3/iBn5iR+3Kpi4aI5FZj6h03FzoR4iIh6YZMuDwJbiKpWEtOIJ+mHmt5+/K/Ef
XNtXfgPwNEMJtiElmdSFFtUEEWCE0lEN38R+79OjXU69BJxpqbky/sbTaqtpIuu2
FLYQY8+ggoMLvZALQvqdwvdpvTAnTo9tSY086MyPvNqdvlMuJse+srTysFVTUejM
vUgtD3hCI9OIcggdev5B2P+VrCBDKPjb6Ua2GAXXniMzt6zcHCPWcys3dddhBhZf
tN3QpMyccQ/O94zhHW2XDC1JJRSunVupZqes6AbMrGniA5JaVsJTwugl9Uiyb+ba
MNcdU9TSTzD1udW6I0HVWVzxygvTncMFXlUe5jaCYWlRazhfxw5XkFfc4Hl4HOIZ
LEwXrRqV+gads/HJQPNrvTK/hyNXHswfi11618Hk6Xa9kQpe2eBJAgFFDSgiwWh+
bWbBduUHwPtFJwDuZEabnPueLJb+uIa95H8b5/mjyYObsfCkIsR3v3zXSLK426sE
ukuuCmiLBWrdRFbHFysMl+/OXLVGYz5FtgSl2LMY85FlFezwjrp05OsmSLz36WWa
NBxiJme23zWhOhTHH6HRhg9YjtazT74/35Pe9LSCpdvy44cbaz3mdyUWs2damOXq
qTxK6jv53jPP2ngDQPrAX0VG74cJ+a6vWJ0OL1djVjJWirj53Gra4/bMZ5X2n0Ot
4/73z+vI6x6qsuKS0vWO+w4yb+cJLufyqWEEzuaS6YmLDDbJ1SISi3d7nvrkngMr
oGXlBuD4ZQcdjHsmi6crmfI+A9Om1tvFg1gb6XmLy4i50qp/J8r7uBGNbMB+wINZ
6KyxA9B/XhG8ALGLowcqWnDwV+w1TNZhi0BjGtDsNq56NvLyZLKNgK6dmF+24nax
BqHR2sKYA3DDfwHDOCw7kTYxNxM3Cs3x+xcpuuuDHmSwB+HA0iNn9/wofmW6AIYN
4QG04OocLY5lOqMDUQS+iQSidDELBPpShBa99taWRWLdzA+jmGl4PqI5rrJGVc62
/X5RdnZdQ8TSXK2jzNKtiBgTlUyb7aIoONckwPPD4ugkqlzoJG39xs1ipdDpzBZH
LmAZvc3M15N6TdeuCP9F8yiT3OSuI1/vZC/0R5F5a+du9yCeLXEW7s2pdX9RFYSM
A4GyEiLeIM/tciKN3HYiOSJzJIrAkEJ169PVUfVVN2NkYVOH8PyPde+E+lAInQDg
imrPCa/KWtiMXjgKKh9Ii3V3YM3juuo/JW/wVbHHDDXFi6KtFa/hNbE9pH6wB8H1
zv2F5rymW1uwJ88YRCLoRdLPvEtkW1wDhG9FnYGWajgiKgEd5uyXT9NKp/uCURLf
Q9Rol6XHNpRZMR4Q/Wf1pcm1v68Qa+x/kl2PfpCn69NSdsjRnKorCYIKgAIeJ6V+
RMovJ8LJdlXKIb7/nNdrxoEaycLDOo80yRLMM0Wc1m/j5yZjxWH/5s0kti1KgO6W
51L1dWi1BHU6W9I6cXtRRQJ3LUEJx1VLvLhd3gqAfjASEkz90DB3SXZmUGISWFUU
i7sb2CYD12GtdFdGdE7hpKTJQDKj6g54lNVFiJXuBPDRwg8HBcGmrLs6Zb5gXi6x
GNoDEbJ+HE07pn2F/4K6BLkRiRTwh1ceuu+E8gxWe81X02vVp8Rh8Re7Wj/iFIAA
2OsvoRkG1Wbn+q3qghyj9WcdVPPtSTA8ViY+xCJ9PvlIuDpill1TCgpJDnX7yuHY
W3Pbp6XgLkNQVCQvwGIAJO/XkSGKVXakitqAAJo9pzC3auUpCJiKl7PIhzfNHw0E
Mmdui1uQ4BQ8cuxYZg0it+qovi/Ec2o0ww+/iwla+eeji0NQ7Fsp/S8H0kvWj9cn
7oehsi9g1t8fx7ifviA4Wyi1H4YeZCsK0gQVsIuCwpZFAwq9Tw7vtlhR0bFqMriq
FYPSvz/hxzYCDRoYygpDKmv2NsFmdM4fIJD9PAQwBEhY7oVYPXJhbYfqqaTzxAEg
cu+hdG9bBk8RRtJiSmpSsK14UUE+/pJOv1T4JeNF1eKD2UVmpJnXNIgIKxHJGDd+
ZuIFQ6kwGKvb8nAkrI+WgwVJyEEgEHsS5oRhbx5gq0UWRE4jVvRcHWTLN/aMUK4/
OCqeyq/Hxx98yAQCCf59cxXEYRWgsCeYS7FmSa240dGP74I2e5B58881CBnp4tJP
oacotqypuPjOsNow8bpLGpLQpPFt3UHRkdBRNirnM4cq6h7vkU6N3l0HLzs+1T0c
ZGY28xAjeyhS3BAZIspgICT/+slBXhM9QslR65NpQigR6iSh7cMNJQl2COkWK2tc
1B7Buoiq5rEnq5PH8SUw4d6LjvHzHaeD5iKFNtBlQX/QBxcc2vj8PBOPu7KCH/vU
jHBqnG45k2ZhAYow97+DV/DZ5CFpbSObEHTdQ/M48JqwCw5QpJNGQEDaB97N/vt2
AFv9ca4yb/H5sd9tKmJJS2FqzLLgIyxUdJaFN8Ah8u45wXitwagQjylfPqdlIZAX
KMyVZYyc3R7pThMp1mMq5qYxdG7UCxC7SMMyeIQYsB0GCOQ7yT2k6n4qnOA3LOlN
sVccRKp4o49ATh4Smg/ZkaCSwqcHBxftW0rW7UJ47kXf2cSdsdZ3qkKTC4GA5+4W
q9T6M5XztdGLsVQDB04MU91KVm7ztbURKR8//HHXOQWDMhCIbJwX4QBEa8kqyVcc
x0NR4yK/PzeTJ2TIkFWcgk6RFK+Q6fcht9EkGUY3p5oogwkgFqYlM3RusjelHJCj
AxbJcB+uY6iiix+RAo65o+ecE5x9R7HiVxzO/AuII6rEWVdZEzB/+OjO3IfjUvIy
fFJT/gR+Wt29XoxRNdA1fJdX8fWBPWOcPDClZ7+EA7y6e3uYcgY0S8Ay5UiPI6S5
N06ZBt9XDz5qzHSy4ZsRRVXZoIzZvMBVr+W+PzOmPDu4yB+CCxlK18I7GBAdDS6b
ECGj5v0rY8MHusKk4byS/SnwHmre0A1/K5ve4WQbzi9BbGabg47bP4RVQmiSGBN4
kku0siv86EHcoMejXIYYUfLz7vfSXCdfuWyCCQN4/HsIt/pQYIhqQIouwEzDDH7T
94iDNXXwxpCJLAU707hLbxbjB8QHMwQkzdXes5KmUQ7lN05JaSvD5bWJEnOmyGfF
OKTIt30FC1dUhZL23GuH5ocSn0Iugazup9YQ9EYrEB5CLyIZGqd25yfeP1mc0l23
mTEwlKr3AxHd4i1MncHxw1dvLuP/bHgxOu30nCBKtbKf2fLYXsxGQqUpR6S53fMZ
b2k1OtfpH/SlS/+zQjNPWDDBZsGALSRBI91r96yIUsSg1UyidhzRD/4S+p0Oi2UZ
g483ESs/9NBO4T1xHAhgwyhuOrJbNVv3QZRQeXwWyvZ+30KSRDYJCSeeRG0/OfGL
uqq9z9EYmd9lxBAw1/fTC4MjKl00114nwtWgE+1c0E/5/0M52ikWEcH9i0OuezPJ
G0MTBQr5QW39tP8x+iOG34R3Tbkj0sJTKQAL2Cf5HNscTVvFSmf7QSJN724YBvSO
yKfHdPNe/TnD9kofcQOBj0FzXt0cO8/H2jUm9+9iidJNXD3AWmhR2YQK8sjUE7RY
muYwUhQ6ITVJVqXpQyYRyGkSJThnyjpFqpAg4JVNwL6wCM7X8hy93HtCb4B3tt71
mcPLDsvXysPELEFLFpW+ZsEiRJvtRLTo0uvkEUHaXIu5DqkprbRUlAsi3BuoE6f0
/yMCfQgcN/E9XFZ6NK67qe7ORB6SWnqnaVxx5TfW0id3/j+z35gZTfleyP2+gEu1
yvpXdAUkPm2xWYRysP4C5fkk0/RzWRgovrydtCm3G9gtBH2QjHYkAdjMqanrIC19
2erH07yBpwLOCHADfCOrB8b2x5nsdoCeehijw19Ad05EcWAgI+GGw1QAoa1+p+xw
B+M3Ahe0eNKaAWgXF7erVluzm3heVhehfurSxs3yPtIL0EH4bmvqr5DCrbi1GJTn
a+YPdAg4N4tJB41pDVvIrQ+ol+poF7e4asy1phmJ3UyBIKJQrIOXMXpbJUnDcU1F
lQGPIWJ+pZUlbgdjgWEjUQxpaLPpMMQbOvUfF+2754lmwT1//M+kmhfRa0jCrd5J
v6LSkkZ7iJ7Gs+SAxa9aIw8mhgd8GmANKVEeEBPLXCOnhAFmnU9e8Ob6lkEeoVP5
MNalTIPJW1tLsOMSOzn3S2+LVpdS57NVXSMjdvTmUcuArDCuGvZSh4Qdn3Nkg6ea
xed0KTGXddizEGj8v9mCvNOV7HlWMxmNLImL7oMzL3fdKzX64mafdqCM2ETYXPVU
aHljpOoBK62UiR1a+fEmqZBNmzPFoxEMt9HhLh9gXUaTDq+2gLW+i4BfeO7uawaw
CxYb0XNK0+ZL4rGqdznrqsFGV2Zmv5cxJNP1dHtFxUrRh6Y4m7xpCVW9EfhX4nOV
VdMSFM4crhQtHsb62/sWlIoJ75cP8SVi+iIAOacOy6H5lFlM6GZ4tvPK4GyeniXx
QUodCAkML9Jxg+mqAKHHdohCCFmsDY3Qi3s15UjK6EP21fqz0lML/sY5x1I2/FUX
FVgjZ3lJ9ka1QjHog8YKAxofxXwfFA3QlxQcYQ6c+AI=
//pragma protect end_data_block
//pragma protect digest_block
EuUUKLOQ9hnFzefQ+VMlHxHo80E=
//pragma protect end_digest_block
//pragma protect end_protected
