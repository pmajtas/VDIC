/******************************************************************************
 * (C) Copyright 2022 AGH UST All Rights Reserved
 ******************************************************************************
 * MODULE NAME: vdic_dut_2022
 * VERSION:     1.3
 * DATE:        24-11-2022
 *
 * ABSTRACT:   DUT module for VDIC 2022 labs.
 *              The DUT is RPN calculator type. The arguments are sent first,
 *              than the operator/command.
 *******************************************************************************
 * HISTORY:
 * 20-10-2022 v1.0 Initial version
 * 03-11-2022 v1.1 Added remaining commands
 * 10-11-2022 v1.2 Modifications:
 *            - corrected bug: zero returned for invalid command
 *            - corrected spec: CMD_AND description
 * 24-11-2022 v1.3 Modifications:
 *            - corrected operation for 10 args
 *            - implemented data parity checking
 * 
 *******************************************************************************
 * INPUTS
 *    clk      - posedge active clock, always running
 *    rst_n    - synchronous reset active low
 *    din      - serial data input
 *    enable_n - chip enable, active low;

 * OUTPUTS
 *    dout       - serial data output
 *    dout_valid - valid flag for serial data output, active high
 *
 *******************************************************************************

 The clock is always active.
 The DUT operates on the posedge of the clock.
 The DUT receives the data when enable_n is active.
 IMPORTANT: din and dout can operate in parallel - DUT has some internal buffering
 implemented.

 --------------------------------------------------------------------------------
 --- Input data
 --------------------------------------------------------------------------------

 The input data is send serially in WORDs.

 The WORD is always 10 bit long. MSB is sent first.
 The WORD sent to the DUT is either DATA type or CONTROL type.

 DATA = 0bbbbbbbbp
 where:
 - b = 0 or 1, PAYLOAD bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 CONTROL = 1bbbbbbbbp
 where:
 - b = 0 or 1, COMMAND bit, total 8 bits, MSB first
 - p = 0 or 1, even parity bit for the 9 bits (total number of 1's in the
 10-bits should be even)

 The COMMAND can be:
 00000000 - CMD_NOP, do nothing, remove the data (reset data stack)
 00000001 - CMD_AND, logic AND of the arguments
 00000010 - CMD_OR, logic OR of the arguments
 00000011 - CMD_XOR, logic XOR of the arguments
 00010000 - CMD_ADD, add the arguments
 00100000 - CMD_SUB, subtract other arguments from the first one

 --------------------------------------------------------------------------------
 --- Output data
 --------------------------------------------------------------------------------

 The DUT responds to each CONTROL word, sending 3 WORDS:
 STATUS, DATA, DATA

 STATUS = 1bbbbbbbbp
 where bbbbbbbb is one of:

 00000000 - S_NO_ERROR - data correctly processed
 00000001 - S_MISSING_DATA - missing input data
 00000010 - S_DATA_STACK_OVERFLOW - maximum number of arguments exceeded
 00000100 - S_OUTPUT_FIFO_OVERFLOW - result dropped not possible to process
 00100000 - S_DATA_PARITY_ERROR - input data or command parity error
 01000000 - S_COMMAND_PARITY_ERROR - input data or command parity error
 10000000 - S_INVALID_COMMAND - unknown command detected

 DATA is defined as in the input.
 PAYLOAD of the DATA is 00000000 if the data was NOT processed correctly.

 *******************************************************************************
 * IMPLEMENTATION STATUS
 *******************************************************************************
 *  <Feature>                        <Is implemented>
 *    command CMD_NOP                   YES
 *    command CMD_AND                   YES
 *    command CMD_OR                    YES
 *    command CMD_XOR                   YES
 *    command CMD_ADD                   YES
 *    command CMD_SUB                   YES
 *    status S_NO_ERROR                 YES
 *    status S_MISSING_DATA              NO
 *    status S_DATA_STACK_OVERFLOW       NO
 *    status S_OUTPUT_FIFO_OVERFLOW      NO
 *    status S_DATA_PARITY_ERROR        YES
 *    status S_COMMAND_PARITY_ERROR      NO
 *    status S_INVALID_COMMAND          YES
 *******************************************************************************
 */

module vdic_dut_2022(clk, rst_n, enable_n, din, dout, dout_valid);
  input clk, rst_n, enable_n, din;
  output dout, dout_valid;
  wire clk, rst_n, enable_n, din;
  wire dout, dout_valid;
  wire [9:0] data_parity_mem;
  wire [7:0] \data_stack_mem[0] ;
  wire [7:0] \data_stack_mem[1] ;
  wire [7:0] \data_stack_mem[2] ;
  wire [7:0] \data_stack_mem[3] ;
  wire [7:0] \data_stack_mem[4] ;
  wire [7:0] \data_stack_mem[5] ;
  wire [7:0] \data_stack_mem[6] ;
  wire [7:0] \data_stack_mem[7] ;
  wire [7:0] \data_stack_mem[8] ;
  wire [7:0] \data_stack_mem[9] ;
  wire [4:0] data_stack_pointer;
  wire [9:0] sh_reg_in;
  wire [4:0] sh_reg_out_bit_counter;
  wire [3:0] sh_bit_cnt;
  wire [2:0] out_fifo_read_pointer;
  wire [9:0] \out_fifo[2][1] ;
  wire [9:0] \out_fifo[1][1] ;
  wire [9:0] \out_fifo[7][1] ;
  wire [9:0] \out_fifo[1][0] ;
  wire [9:0] \out_fifo[4][0] ;
  wire [9:0] \out_fifo[2][0] ;
  wire [9:0] \out_fifo[0][0] ;
  wire [9:0] \out_fifo[6][0] ;
  wire [9:0] \out_fifo[3][0] ;
  wire [9:0] \out_fifo[5][0] ;
  wire [9:0] \out_fifo[7][0] ;
  wire [9:0] \out_fifo[0][1] ;
  wire [9:0] \out_fifo[3][1] ;
  wire [9:0] \out_fifo[5][1] ;
  wire [9:0] \out_fifo[7][2] ;
  wire [9:0] \out_fifo[5][2] ;
  wire [9:0] \out_fifo[3][2] ;
  wire [9:0] \out_fifo[6][2] ;
  wire [9:0] \out_fifo[0][2] ;
  wire [9:0] \out_fifo[6][1] ;
  wire [9:0] \out_fifo[2][2] ;
  wire [9:0] \out_fifo[4][2] ;
  wire [9:0] \out_fifo[1][2] ;
  wire [9:0] \out_fifo[4][1] ;
  wire [2:0] out_fifo_write_pointer;
  wire [29:0] sh_reg_out;
  wire n_16065, n_16066, n_16067, n_16068, n_16069, n_16074, n_16075,
       n_16076;
  wire n_16077, n_16078, n_16079, n_16080, n_16081, n_16082, n_16083,
       n_16084;
  wire n_16085, n_16086, n_16087, n_16088, n_16089, n_16090, n_16091,
       n_16092;
  wire n_16093, n_16094, n_16095, n_16099, n_16100, n_16103, n_16105,
       n_16106;
  wire n_16107, n_16108, n_16109, n_16110, n_16111, n_16112, n_16113,
       n_16114;
  wire n_16115, n_16116, n_16117, n_16118, n_16119, n_16120, n_16121,
       n_16122;
  wire n_16123, n_16124, n_16125, n_16126, n_16127, n_16128, n_16129,
       n_16130;
  wire n_16131, n_16132, n_16133, n_16134, n_16135, n_16136, n_16137,
       n_16139;
  wire n_16140, n_16141, n_16142, n_16143, n_16144, n_16145, n_16146,
       n_16147;
  wire n_16148, n_16149, n_16150, n_16151, n_16152, n_16153, n_16154,
       n_16155;
  wire n_16156, n_16157, n_16158, n_16159, n_16160, n_16161, n_16162,
       n_16163;
  wire n_16164, n_16165, n_16166, n_16167, n_16168, n_16169, n_16170,
       n_16171;
  wire n_16172, n_16173, n_16174, n_16175, n_16176, n_16177, n_16178,
       n_16179;
  wire n_16180, n_16181, n_16182, n_16183, n_16184, n_16185, n_16186,
       n_16187;
  wire n_16188, n_16189, n_16190, n_16191, n_16192, n_16193, n_16194,
       n_16195;
  wire n_16196, n_16197, n_16198, n_16199, n_16200, n_16201, n_16202,
       n_16203;
  wire n_16204, n_16205, n_16206, n_16207, n_16208, n_16209, n_16210,
       n_16211;
  wire n_16212, n_16213, n_16214, n_16215, n_16216, n_16217, n_16218,
       n_16219;
  wire n_16220, n_16221, n_16222, n_16223, n_16224, n_16225, n_16226,
       n_16227;
  wire n_16228, n_16229, n_16230, n_16231, n_16232, n_16233, n_16234,
       n_16235;
  wire n_16236, n_16237, n_16238, n_16239, n_16240, n_16241, n_16242,
       n_16243;
  wire n_16244, n_16245, n_16246, n_16247, n_16248, n_16249, n_16250,
       n_16251;
  wire n_16252, n_16253, n_16254, n_16255, n_16256, n_16257, n_16258,
       n_16259;
  wire n_16260, n_16261, n_16262, n_16263, n_16264, n_16265, n_16266,
       n_16267;
  wire n_16268, n_16269, n_16270, n_16271, n_16272, n_16273, n_16274,
       n_16275;
  wire n_16276, n_16277, n_16278, n_16279, n_16280, n_16281, n_16282,
       n_16283;
  wire n_16284, n_16285, n_16286, n_16287, n_16288, n_16289, n_16290,
       n_16291;
  wire n_16292, n_16293, n_16294, n_16295, n_16296, n_16297, n_16298,
       n_16299;
  wire n_16300, n_16301, n_16302, n_16303, n_16304, n_16305, n_16306,
       n_16307;
  wire n_16308, n_16309, n_16310, n_16311, n_16312, n_16313, n_16314,
       n_16315;
  wire n_16316, n_16317, n_16318, n_16319, n_16320, n_16321, n_16322,
       n_16323;
  wire n_16324, n_16325, n_16326, n_16327, n_16328, n_16329, n_16330,
       n_16331;
  wire n_16332, n_16333, n_16334, n_16335, n_16336, n_16337, n_16338,
       n_16339;
  wire n_16340, n_16341, n_16342, n_16343, n_16344, n_16345, n_16346,
       n_16347;
  wire n_16348, n_16349, n_16350, n_16351, n_16352, n_16353, n_16354,
       n_16355;
  wire n_16356, n_16357, n_16358, n_16359, n_16360, n_16361, n_16362,
       n_16363;
  wire n_16364, n_16365, n_16366, n_16367, n_16368, n_16369, n_16370,
       n_16371;
  wire n_16372, n_16373, n_16374, n_16375, n_16376, n_16377, n_16378,
       n_16379;
  wire n_16380, n_16381, n_16382, n_16383, n_16384, n_16385, n_16386,
       n_16387;
  wire n_16388, n_16389, n_16390, n_16391, n_16392, n_16393, n_16394,
       n_16395;
  wire n_16396, n_16397, n_16398, n_16399, n_16400, n_16401, n_16402,
       n_16403;
  wire n_16404, n_16405, n_16406, n_16407, n_16408, n_16409, n_16410,
       n_16411;
  wire n_16412, n_16413, n_16414, n_16415, n_16416, n_16417, n_16418,
       n_16419;
  wire n_16420, n_16421, n_16422, n_16423, n_16424, n_16425, n_16426,
       n_16427;
  wire n_16428, n_16429, n_16430, n_16431, n_16432, n_16433, n_16434,
       n_16435;
  wire n_16436, n_16437, n_16438, n_16439, n_16440, n_16441, n_16442,
       n_16443;
  wire n_16444, n_16445, n_16446, n_16447, n_16448, n_16449, n_16450,
       n_16451;
  wire n_16452, n_16453, n_16454, n_16455, n_16456, n_16457, n_16458,
       n_16459;
  wire n_16460, n_16461, n_16462, n_16463, n_16464, n_16465, n_16466,
       n_16467;
  wire n_16468, n_16469, n_16470, n_16471, n_16472, n_16473, n_16474,
       n_16475;
  wire n_16476, n_16477, n_16478, n_16479, n_16480, n_16481, n_16482,
       n_16483;
  wire n_16484, n_16485, n_16486, n_16487, n_16488, n_16489, n_16490,
       n_16491;
  wire n_16492, n_16493, n_16494, n_16495, n_16496, n_16497, n_16498,
       n_16499;
  wire n_16500, n_16501, n_16502, n_16503, n_16504, n_16505, n_16506,
       n_16507;
  wire n_16508, n_16509, n_16510, n_16511, n_16512, n_16513, n_16514,
       n_16515;
  wire n_16516, n_16517, n_16518, n_16519, n_16520, n_16521, n_16522,
       n_16523;
  wire n_16524, n_16525, n_16526, n_16527, n_16528, n_16529, n_16530,
       n_16531;
  wire n_16532, n_16533, n_16535, n_16536, n_16537, n_16538, n_16539,
       n_16540;
  wire n_16541, n_16542, n_16543, n_16544, n_16545, n_16546, n_16547,
       n_16548;
  wire n_16549, n_16550, n_16551, n_16552, n_16553, n_16554, n_16555,
       n_16556;
  wire n_16557, n_16558, n_16559, n_16560, n_16561, n_16562, n_16563,
       n_16564;
  wire n_16565, n_16566, n_16567, n_16568, n_16569, n_16570, n_16571,
       n_16572;
  wire n_16573, n_16574, n_16575, n_16576, n_16577, n_16578, n_16579,
       n_16580;
  wire n_16581, n_16582, n_16583, n_16584, n_16585, n_16586, n_16587,
       n_16588;
  wire n_16589, n_16590, n_16591, n_16592, n_16593, n_16594, n_16595,
       n_16596;
  wire n_16597, n_16598, n_16599, n_16600, n_16601, n_16602, n_16603,
       n_16604;
  wire n_16605, n_16606, n_16607, n_16608, n_16609, n_16610, n_16611,
       n_16612;
  wire n_16613, n_16614, n_16615, n_16616, n_16617, n_16618, n_16619,
       n_16620;
  wire n_16621, n_16622, n_16623, n_16624, n_16625, n_16626, n_16627,
       n_16628;
  wire n_16629, n_16630, n_16631, n_16632, n_16633, n_16634, n_16635,
       n_16636;
  wire n_16637, n_16638, n_16639, n_16640, n_16641, n_16642, n_16643,
       n_16644;
  wire n_16645, n_16646, n_16647, n_16648, n_16649, n_16650, n_16651,
       n_16652;
  wire n_16653, n_16654, n_16655, n_16656, n_16657, n_16658, n_16659,
       n_16660;
  wire n_16661, n_16662, n_16663, n_16664, n_16665, n_16666, n_16667,
       n_16668;
  wire n_16669, n_16670, n_16671, n_16672, n_16673, n_16674, n_16675,
       n_16676;
  wire n_16677, n_16678, n_16679, n_16680, n_16681, n_16682, n_16683,
       n_16684;
  wire n_16685, n_16686, n_16687, n_16688, n_16689, n_16690, n_16691,
       n_16692;
  wire n_16693, n_16694, n_16695, n_16696, n_16697, n_16698, n_16699,
       n_16700;
  wire n_16701, n_16702, n_16703, n_16704, n_16705, n_16706, n_16707,
       n_16708;
  wire n_16709, n_16710, n_16711, n_16712, n_16713, n_16714, n_16715,
       n_16716;
  wire n_16717, n_16718, n_16719, n_16720, n_16721, n_16722, n_16723,
       n_16724;
  wire n_16725, n_16726, n_16727, n_16728, n_16729, n_16730, n_16731,
       n_16732;
  wire n_16733, n_16734, n_16735, n_16736, n_16737, n_16738, n_16739,
       n_16740;
  wire n_16741, n_16742, n_16743, n_16744, n_16745, n_16746, n_16747,
       n_16748;
  wire n_16749, n_16750, n_16751, n_16752, n_16753, n_16754, n_16755,
       n_16756;
  wire n_16757, n_16758, n_16760, n_16761, n_16762, n_16763, n_16764,
       n_16765;
  wire n_16766, n_16767, n_16768, n_16769, n_16770, n_16771, n_16772,
       n_16773;
  wire n_16774, n_16775, n_16776, n_16777, n_16778, n_16779, n_16780,
       n_16781;
  wire n_16782, n_16783, n_16784, n_16785, n_16786, n_16787, n_16788,
       n_16789;
  wire n_16790, n_16791, n_16792, n_16793, n_16794, n_16795, n_16796,
       n_16797;
  wire n_16798, n_16799, n_16800, n_16801, n_16802, n_16803, n_16804,
       n_16805;
  wire n_16806, n_16807, n_16808, n_16809, n_16810, n_16811, n_16812,
       n_16813;
  wire n_16814, n_16815, n_16816, n_16817, n_16818, n_16819, n_16820,
       n_16821;
  wire n_16822, n_16823, n_16824, n_16825, n_16826, n_16827, n_16828,
       n_16829;
  wire n_16830, n_16831, n_16832, n_16833, n_16834, n_16835, n_16836,
       n_16837;
  wire n_16838, n_16839, n_16840, n_16841, n_16842, n_16843, n_16844,
       n_16845;
  wire n_16846, n_16847, n_16848, n_16849, n_16850, n_16851, n_16852,
       n_16853;
  wire n_16854, n_16855, n_16856, n_16857, n_16858, n_16859, n_16860,
       n_16861;
  wire n_16862, n_16863, n_16864, n_16865, n_16866, n_16867, n_16868,
       n_16869;
  wire n_16870, n_16871, n_16872, n_16873, n_16874, n_16875, n_16876,
       n_16877;
  wire n_16878, n_16879, n_16880, n_16881, n_16882, n_16883, n_16889,
       n_16890;
  wire n_16891, n_16892, n_16893, n_16894, n_16895, n_16896, n_16897,
       n_16898;
  wire n_16899, n_16900, n_16901, n_16902, n_16903, n_16904, n_16905,
       n_16906;
  wire n_16907, n_16908, n_16909, n_16910, n_16911, n_16912, n_16913,
       n_16914;
  wire n_16915, n_16916, n_16917, n_16918, n_16919, n_16920, n_16921,
       n_16922;
  wire n_16923, n_16924, n_16925, n_16926, n_16927, n_16928, n_16929,
       n_16930;
  wire n_16931, n_16932, n_16933, n_16934, n_16935, n_16936, n_16937,
       n_16938;
  wire n_16939, n_16940, n_16941, n_16942, n_16943, n_16944, n_16945,
       n_16946;
  wire n_16947, n_16948, n_16949, n_16950, n_16951, n_16952, n_16953,
       n_16954;
  wire n_16955, n_16956, n_16957, n_16958, n_16959, n_16960, n_16961,
       n_16962;
  wire n_16963, n_16964, n_16965, n_16966, n_16967, n_16968, n_16969,
       n_16970;
  wire n_16971, n_16972, n_16973, n_16974, n_16975, n_16976, n_16977,
       n_16978;
  wire n_16979, n_16980, n_16981, n_16982, n_16983, n_16984, n_16985,
       n_16986;
  wire n_16987, n_16988, n_16989, n_16990, n_16991, n_16992, n_16993,
       n_16994;
  wire n_16995, n_16996, n_16997, n_16998, n_16999, n_17000, n_17001,
       n_17002;
  wire n_17003, n_17004, n_17005, n_17006, n_17007, n_17008, n_17009,
       n_17010;
  wire n_17011, n_17012, n_17013, n_17014, n_17015, n_17016, n_17017,
       n_17018;
  wire n_17019, n_17020, n_17021, n_17022, n_17023, n_17024, n_17025,
       n_17026;
  wire n_17027, n_17028, n_17029, n_17030, n_17031, n_17032, n_17033,
       n_17034;
  wire n_17035, n_17036, n_17037, n_17038, n_17039, n_17040, n_17041,
       n_17042;
  wire n_17043, n_17044, n_17045, n_17046, n_17047, n_17048, n_17049,
       n_17050;
  wire n_17051, n_17052, n_17053, n_17055, n_17056, n_17057, n_17058,
       n_17059;
  wire n_17060, n_17061, n_17063, n_17064, n_17065, n_17066, n_17067,
       n_17068;
  wire n_17069, n_17070, n_17071, n_17072, n_17073, n_17074, n_17075,
       n_17076;
  wire n_17077, n_17078, n_17079, n_17080, n_17081, n_17082, n_17083,
       n_17084;
  wire n_17085, n_17086, n_17087, n_17088, n_17089, n_17090, n_17091,
       n_17092;
  wire n_17093, n_17094, n_17095, n_17096, n_17097, n_17098, n_17099,
       n_17100;
  wire n_17101, n_17102, n_17103, n_17104, n_17105, n_17106, n_17107,
       n_17108;
  wire n_17109, n_17110, n_17111, n_17112, n_17113, n_17114, n_17115,
       n_17116;
  wire n_17117, n_17118, n_17119, n_17120, n_17121, n_17125, n_17126,
       n_17127;
  wire n_17128, n_17129, n_17130, n_17131, n_17132, n_17133, n_17134,
       n_17135;
  wire n_17136, n_17137, n_17138, n_17139, n_17140, n_17141, n_17142,
       n_17143;
  wire n_17144, n_17145, n_17146, n_17147, n_17245, n_17260, n_17265,
       n_17284;
  wire n_17286, n_17287, n_17290, n_17293, n_17294, n_17296, n_17298,
       n_17300;
  wire n_17303, n_17310, n_17315, n_17316, n_17317, n_17318, n_17319,
       n_17320;
  wire n_17321, n_17322, n_17323, n_17324, n_17325, n_17326, n_17327,
       n_17328;
  wire n_17329, n_17330, n_17331, n_17332, n_17333, n_17334, n_17335,
       n_17336;
  wire n_17337, n_17338, n_17339, n_17340, n_17341, n_17342, n_17343,
       n_17344;
  wire n_17345, n_17346, n_17347, n_17348, n_17349, n_17350, n_17351,
       n_17352;
  wire n_17353, n_17354, n_17355, n_17356, n_17357, n_17358, n_17359,
       n_17360;
  wire n_17361, n_17362, n_17363, n_17364, n_17365, n_17366, n_17369,
       n_17370;
  wire n_17371, n_17372, n_17373, n_17374, n_17375, n_17376, n_17377,
       n_17378;
  wire n_17379, n_17380, n_17381, n_17382, n_17383, n_17384, n_17385,
       n_17386;
  wire n_17387, n_17388, n_17389, n_17390, n_17391, n_17392, n_17393,
       n_17394;
  wire n_17395, n_17396, n_17397, n_17398, n_17399, n_17400, n_17402,
       n_17403;
  wire n_17404, n_17405, n_17406, n_17407, n_17408, n_17409, n_17410,
       n_17411;
  wire n_17412, n_17413, n_17414, n_17415, n_17416, n_17417, n_17418,
       n_17419;
  wire n_17421, n_17422, n_17423, n_17424, n_17425, n_17426, n_17427,
       n_17429;
  wire n_17430, n_17431, n_17432, n_17433, n_17435, n_17436, n_17437,
       n_17438;
  wire n_17439, n_17440, n_17441, n_17442, n_17443, n_17444, n_17445,
       n_17446;
  wire n_17447, n_17448, n_17449, n_17450, n_17452, n_17453, n_17454,
       n_17456;
  wire n_17457, n_17459, n_17460, n_17461, n_17462, n_17464, n_17465,
       n_17466;
  wire n_17467, n_17481, n_17501, n_17507, n_17508, n_17510, n_17511,
       n_17512;
  wire n_17634, n_17635, n_17636, n_17638, n_17640, n_17642, n_17643,
       n_17644;
  wire n_17645, n_17646, n_17647, n_17650, n_17651, n_17653, n_17654,
       n_17655;
  wire n_17657, n_17658, n_17660, n_17662, n_17664, n_17665, n_17667,
       n_17668;
  wire n_17669, n_17671, n_17672, n_17674, n_17676, n_17678, n_17680,
       n_17682;
  wire n_17684, n_17686, n_17687, n_17689, n_17690, n_17691, n_17693,
       n_17694;
  wire n_17695, n_17696, n_17697, n_17698, n_17699, n_17700, n_17701,
       n_17702;
  wire n_17703, n_17704, n_17705, n_17706, n_17707, n_17708, n_17710,
       n_17711;
  wire n_17713, n_17714, n_17715, n_17716, n_17717, n_17718, n_17719,
       n_17720;
  wire n_17722, n_17723, n_17724, n_17725, n_17726, n_17727, n_17728,
       n_17729;
  wire n_17730, n_17731, n_17732, n_17733, n_17734, n_17735, n_17736,
       n_17737;
  wire n_17738, n_17739, n_17740, n_17741, n_17742, n_17743, n_17744,
       n_17745;
  wire n_17746, n_17747, n_17748, n_17749, n_17750, n_17751, n_17752,
       n_17753;
  wire n_17754, n_17755, n_17756, n_17757, n_17758, n_17759, n_17760,
       n_17761;
  wire n_17762, n_17763, n_17771, n_17772, n_17799, n_17800, n_17801,
       n_17802;
  wire n_17803, n_17804, n_17805, n_17806, n_17816, n_17817, n_17818,
       n_17823;
  wire n_17824, n_17841, n_17842, n_17843, n_17844, n_17845, n_17846,
       n_17847;
  wire n_17848, n_17851, n_17858, n_17859, n_17860, n_17863, n_17870,
       n_17871;
  wire n_17872, n_17883, n_17884, n_17889, n_17890, n_17893, n_17896,
       n_17899;
  wire n_17902, n_17905, n_17908, n_17911, n_17916, n_17917, n_17922,
       n_17923;
  wire n_17926, n_17929, n_17932, n_17935, n_17942, n_17943, n_17944,
       n_17949;
  wire n_17950, n_17953, n_17956, n_17963, n_17964, n_17965, n_17970,
       n_17971;
  wire n_17974, n_17977, n_17980, n_17985, n_17986, n_18019, n_18020,
       n_18021;
  wire n_18022, n_18023, n_18024, n_18025, n_18026, n_18027, n_18028,
       n_18029;
  wire n_18030, n_18031, n_18032, n_18033, n_18034, n_18037, n_18040,
       n_18043;
  wire n_18046, n_18059, n_18060, n_18061, n_18062, n_18063, n_18064,
       n_18079;
  wire n_18080, n_18081, n_18082, n_18083, n_18084, n_18085, n_18088,
       n_18091;
  wire n_18100, n_18101, n_18103, n_18106, n_18121, n_18122, n_18123,
       n_18124;
  wire n_18125, n_18126, n_18127, n_18142, n_18143, n_18144, n_18145,
       n_18146;
  wire n_18147, n_18148, n_18151, n_18154, n_18159, n_18160, n_18175,
       n_18176;
  wire n_18177, n_18178, n_18179, n_18180, n_18181, n_18196, n_18197,
       n_18198;
  wire n_18199, n_18200, n_18201, n_18202, n_18205, n_18220, n_18221,
       n_18222;
  wire n_18223, n_18224, n_18225, n_18226, n_18241, n_18242, n_18243,
       n_18244;
  wire n_18245, n_18246, n_18247, n_18250, n_18253, n_18262, n_18263,
       n_18264;
  wire n_18265, n_18274, n_18275, n_18276, n_18277, n_18286, n_18287,
       n_18288;
  wire n_18289, n_18298, n_18299, n_18300, n_18301, n_18310, n_18311,
       n_18312;
  wire n_18313, n_18322, n_18323, n_18324, n_18325, n_18335, n_18336,
       n_18337;
  wire n_18346, n_18347, n_18348, n_18349, n_18354, n_18355, n_18358,
       n_18361;
  wire n_18367, n_18370, n_18376, n_18379, n_18382, n_18387, n_18388,
       n_18393;
  wire n_18394, n_18399, n_18400, n_18405, n_18406, n_18411, n_18412,
       n_18417;
  wire n_18418, n_18423, n_18424, n_18429, n_18430, n_18435, n_18436,
       n_18443;
  wire n_18444, n_18445, n_18448, n_18455, n_18456, n_18457, n_18464,
       n_18465;
  wire n_18466, n_18469, n_18472, n_18475, n_18478, n_18481, n_18486,
       n_18487;
  wire n_18512, n_18513, n_18514, n_18515, n_18516, n_18517, n_18518,
       n_18519;
  wire n_18520, n_18521, n_18522, n_18523, n_18526, n_18537, n_18538,
       n_18539;
  wire n_18540, n_18541, n_18546, n_18547, n_18556, n_18557, n_18558,
       n_18559;
  wire n_18566, n_18567, n_18568, n_18571, n_18574, n_18577, n_18580,
       n_18583;
  wire n_18586, n_18591, n_18592, n_18597, n_18598, n_18603, n_18604,
       n_18609;
  wire n_18610, n_18615, n_18616, n_18621, n_18622, n_18627, n_18628,
       n_18633;
  wire n_18634, n_18639, n_18640, n_18645, n_18646, n_18651, n_18652,
       n_18657;
  wire n_18658, n_18663, n_18664, n_18669, n_18670, n_18675, n_18676,
       n_18681;
  wire n_18682, n_18687, n_18688, n_18693, n_18694, n_18699, n_18700,
       n_18705;
  wire n_18706, n_18711, n_18712, n_18717, n_18718, n_18723, n_18724,
       n_18729;
  wire n_18730, n_18735, n_18736, n_18741, n_18742, n_18747, n_18748,
       n_18753;
  wire n_18754, n_18759, n_18760, n_18765, n_18766, n_18771, n_18772,
       n_18777;
  wire n_18778, n_18783, n_18784, n_18789, n_18790, n_18795, n_18796,
       n_18801;
  wire n_18802, n_18807, n_18808, n_18813, n_18814, n_18819, n_18820,
       n_18825;
  wire n_18826, n_18831, n_18832, n_18837, n_18838, n_18843, n_18844,
       n_18849;
  wire n_18850, n_18855, n_18856, n_18861, n_18862, n_18867, n_18868,
       n_18873;
  wire n_18874, n_18879, n_18880, n_18885, n_18886, n_18891, n_18892,
       n_18897;
  wire n_18898, n_18903, n_18904, n_18911, n_18912, n_18913, n_18916,
       n_18919;
  wire n_18940, n_18941, n_18942, n_18943, n_18944, n_18945, n_18946,
       n_18947;
  wire n_18948, n_18949, n_18972, n_18973, n_18974, n_18975, n_18976,
       n_18977;
  wire n_18978, n_18979, n_18980, n_18981, n_18982, n_19003, n_19004,
       n_19005;
  wire n_19006, n_19007, n_19008, n_19009, n_19010, n_19011, n_19012,
       n_19033;
  wire n_19034, n_19035, n_19036, n_19037, n_19038, n_19039, n_19040,
       n_19041;
  wire n_19042, n_19063, n_19064, n_19065, n_19066, n_19067, n_19068,
       n_19069;
  wire n_19070, n_19071, n_19072, n_19093, n_19094, n_19095, n_19096,
       n_19097;
  wire n_19098, n_19099, n_19100, n_19101, n_19102, n_19105, n_19114,
       n_19115;
  wire n_19116, n_19117, n_19126, n_19127, n_19128, n_19129, n_19132,
       n_19135;
  wire n_19142, n_19143, n_19144, n_19147, n_19150, n_19155, n_19156,
       n_19161;
  wire n_19162, n_19167, n_19168, n_19173, n_19174, n_19179, n_19180,
       n_19185;
  wire n_19186, n_19191, n_19192, n_19197, n_19198, n_19203, n_19204,
       n_19209;
  wire n_19210, n_19215, n_19216, n_19221, n_19222, n_19227, n_19228,
       n_19233;
  wire n_19234, n_19239, n_19240, n_19245, n_19246, n_19251, n_19252,
       n_19257;
  wire n_19258, n_19263, n_19264, n_19269, n_19270, n_19275, n_19276,
       n_19281;
  wire n_19282, n_19287, n_19288, n_19293, n_19294, n_19299, n_19300,
       n_19305;
  wire n_19306, n_19311, n_19312, n_19317, n_19318, n_19323, n_19324,
       n_19329;
  wire n_19330, n_19335, n_19336, n_19341, n_19342, n_19347, n_19348,
       n_19353;
  wire n_19354, n_19359, n_19360, n_19365, n_19366, n_19371, n_19372,
       n_19377;
  wire n_19378, n_19383, n_19384, n_19389, n_19390, n_19395, n_19396,
       n_19401;
  wire n_19402, n_19407, n_19408, n_19413, n_19414, n_19419, n_19420,
       n_19425;
  wire n_19435, n_19436, n_19437, n_19438, n_19447, n_19448, n_19449,
       n_19450;
  wire n_19461, n_19462, n_19463, n_19464, n_19465, n_19470, n_19471,
       n_19474;
  wire n_19477, n_19482, n_19483, n_19488, n_19489, n_19494, n_19495,
       n_19500;
  wire n_19501, n_19506, n_19507, n_19512, n_19513, n_19518, n_19519,
       n_19524;
  wire n_19525, n_19530, n_19531, n_19536, n_19537, n_19542, n_19543,
       n_19548;
  wire n_19549, n_19554, n_19555, n_19560, n_19561, n_19566, n_19567,
       n_19572;
  wire n_19573, n_19578, n_19579, n_19584, n_19585, n_19590, n_19591,
       n_19596;
  wire n_19597, n_19626, n_19627, n_19628, n_19629, n_19630, n_19631,
       n_19632;
  wire n_19633, n_19634, n_19635, n_19636, n_19637, n_19638, n_19639,
       n_19672;
  wire n_19673, n_19674, n_19675, n_19676, n_19677, n_19678, n_19679,
       n_19680;
  wire n_19681, n_19682, n_19683, n_19684, n_19685, n_19686, n_19687,
       n_19720;
  wire n_19721, n_19722, n_19723, n_19724, n_19725, n_19726, n_19727,
       n_19728;
  wire n_19729, n_19730, n_19731, n_19732, n_19733, n_19734, n_19735,
       n_19768;
  wire n_19769, n_19770, n_19771, n_19772, n_19773, n_19774, n_19775,
       n_19776;
  wire n_19777, n_19778, n_19779, n_19780, n_19781, n_19782, n_19783,
       n_19816;
  wire n_19817, n_19818, n_19819, n_19820, n_19821, n_19822, n_19823,
       n_19824;
  wire n_19825, n_19826, n_19827, n_19828, n_19829, n_19830, n_19831,
       n_19864;
  wire n_19865, n_19866, n_19867, n_19868, n_19869, n_19870, n_19871,
       n_19872;
  wire n_19873, n_19874, n_19875, n_19876, n_19877, n_19878, n_19879,
       n_19912;
  wire n_19913, n_19914, n_19915, n_19916, n_19917, n_19918, n_19919,
       n_19920;
  wire n_19921, n_19922, n_19923, n_19924, n_19925, n_19926, n_19927,
       n_19960;
  wire n_19961, n_19962, n_19963, n_19964, n_19965, n_19966, n_19967,
       n_19968;
  wire n_19969, n_19970, n_19971, n_19972, n_19973, n_19974, n_19975,
       n_20008;
  wire n_20009, n_20010, n_20011, n_20012, n_20013, n_20014, n_20015,
       n_20016;
  wire n_20017, n_20018, n_20019, n_20020, n_20021, n_20022, n_20023,
       n_20056;
  wire n_20057, n_20058, n_20059, n_20060, n_20061, n_20062, n_20063,
       n_20064;
  wire n_20065, n_20066, n_20067, n_20068, n_20069, n_20070, n_20071,
       n_20104;
  wire n_20105, n_20106, n_20107, n_20108, n_20109, n_20110, n_20111,
       n_20112;
  wire n_20113, n_20114, n_20115, n_20116, n_20117, n_20118, n_20119,
       n_20152;
  wire n_20153, n_20154, n_20155, n_20156, n_20157, n_20158, n_20159,
       n_20160;
  wire n_20161, n_20162, n_20163, n_20164, n_20165, n_20166, n_20167,
       n_20200;
  wire n_20201, n_20202, n_20203, n_20204, n_20205, n_20206, n_20207,
       n_20208;
  wire n_20209, n_20210, n_20211, n_20212, n_20213, n_20214, n_20215,
       n_20248;
  wire n_20249, n_20250, n_20251, n_20252, n_20253, n_20254, n_20255,
       n_20256;
  wire n_20257, n_20258, n_20259, n_20260, n_20261, n_20262, n_20263,
       n_20296;
  wire n_20297, n_20298, n_20299, n_20300, n_20301, n_20302, n_20303,
       n_20304;
  wire n_20305, n_20306, n_20307, n_20308, n_20309, n_20310, n_20311,
       n_20344;
  wire n_20345, n_20346, n_20347, n_20348, n_20349, n_20350, n_20351,
       n_20352;
  wire n_20353, n_20354, n_20355, n_20356, n_20357, n_20358, n_20359,
       n_20392;
  wire n_20393, n_20394, n_20395, n_20396, n_20397, n_20398, n_20399,
       n_20400;
  wire n_20401, n_20402, n_20403, n_20404, n_20405, n_20406, n_20407,
       n_20440;
  wire n_20441, n_20442, n_20443, n_20444, n_20445, n_20446, n_20447,
       n_20448;
  wire n_20449, n_20450, n_20451, n_20452, n_20453, n_20454, n_20455,
       n_20488;
  wire n_20489, n_20490, n_20491, n_20492, n_20493, n_20494, n_20495,
       n_20496;
  wire n_20497, n_20498, n_20499, n_20500, n_20501, n_20502, n_20503,
       n_20536;
  wire n_20537, n_20538, n_20539, n_20540, n_20541, n_20542, n_20543,
       n_20544;
  wire n_20545, n_20546, n_20547, n_20548, n_20549, n_20550, n_20551,
       n_20584;
  wire n_20585, n_20586, n_20587, n_20588, n_20589, n_20590, n_20591,
       n_20592;
  wire n_20593, n_20594, n_20595, n_20596, n_20597, n_20598, n_20599,
       n_20632;
  wire n_20633, n_20634, n_20635, n_20636, n_20637, n_20638, n_20639,
       n_20640;
  wire n_20641, n_20642, n_20643, n_20644, n_20645, n_20646, n_20647,
       n_20680;
  wire n_20681, n_20682, n_20683, n_20684, n_20685, n_20686, n_20687,
       n_20688;
  wire n_20689, n_20690, n_20691, n_20692, n_20693, n_20694, n_20695,
       n_20700;
  wire n_20701, n_20706, n_20707, n_20712, n_20713, n_20718, n_20719,
       n_20724;
  wire n_20725, n_20732, n_20733, n_20734, n_20739, n_20740, n_20745,
       n_20746;
  wire n_20751, n_20752, n_20757, n_20758, n_20763, n_20771, n_20772,
       n_20773;
  wire n_20780, n_20781, n_20782, n_20789, n_20790, n_20791, n_20796,
       n_20797;
  wire n_20802, n_20803, n_20808, n_20809, n_20814, n_20815, n_20820,
       n_20828;
  wire n_20829, n_20830, n_20837, n_20838, n_20839, n_20846, n_20847,
       n_20848;
  wire n_20855, n_20856, n_20857, n_20862, n_20863, n_20868, n_20869,
       n_20874;
  wire n_20875, n_20880, n_20881, n_20886, n_20887, n_20894, n_20895,
       n_20896;
  wire n_20910, n_20918, n_20919, n_20920, n_20925, n_20926, n_20931,
       n_20932;
  wire n_20937, n_20938, n_20943, n_20944, n_20949, n_20950, n_20955,
       n_20956;
  wire n_20961, n_20967, n_20973, n_20974, n_20979, n_20980, n_20985,
       n_20986;
  wire n_20997, n_20998, n_20999, n_21000, n_21001, n_21014, n_21015,
       n_21016;
  wire n_21017, n_21018, n_21019, n_21024, n_21025, n_21030, n_21031,
       n_21036;
  wire n_21037, n_21042, n_21043, n_21048, n_21049, n_21054, n_21055,
       n_21060;
  wire n_21066, n_21072, n_21073, n_21078, n_21079, n_21084, n_21085,
       n_21098;
  wire n_21099, n_21100, n_21101, n_21102, n_21103, n_21108, n_21109,
       n_21112;
  wire n_21117, n_21118, n_21123, n_21124, n_21129, n_21130, n_21135,
       n_21136;
  wire n_21141, n_21142, n_21147, n_21148, n_21153, n_21154, n_21159,
       n_21160;
  wire n_21165, n_21166, n_21171, n_21172, n_21177, n_21178, n_21183,
       n_21184;
  wire n_21191, n_21192, n_21193, n_21198, n_21204, n_21205, n_21212,
       n_21213;
  wire n_21214, n_21219, n_21220, n_21225, n_21226, n_21231, n_21232,
       n_21237;
  wire n_21238, n_21243, n_21247, n_21252, n_21253, n_21260, n_21261,
       n_21262;
  wire n_21267, n_21268, n_21273, n_21274, n_21279, n_21280, n_21285,
       n_21286;
  wire n_21291, n_21292, n_21297, n_21298, n_21303, n_21304, n_21309,
       n_21310;
  wire n_21315, n_21316, n_21321, n_21327, n_21328, n_21331, n_21336,
       n_21337;
  wire n_21340, n_21351, n_21352, n_21353, n_21354, n_21355, n_21360,
       n_21361;
  wire n_21366, n_21367, n_21374, n_21375, n_21376, n_21381, n_21382,
       n_21387;
  wire n_21388, n_21393, n_21394, n_21399, n_21400, n_21405, n_21406,
       n_21411;
  wire n_21412, n_21417, n_21418, n_21423, n_21424, n_21429, n_21430,
       n_21435;
  wire n_21436, n_21441, n_21447, n_21448, n_21451, n_21454, n_21459,
       n_21460;
  wire n_21465, n_21466, n_21471, n_21472, n_21477, n_21478, n_21483,
       n_21484;
  wire n_21489, n_21490, n_21495, n_21496, n_21501, n_21513, n_21514,
       n_21515;
  wire n_21516, n_21517, n_21520, n_21525, n_21526, n_21531, n_21532,
       n_21537;
  wire n_21538, n_21543, n_21544, n_21549, n_21550, n_21555, n_21556,
       n_21563;
  wire n_21564, n_21565, n_21570, n_21571, n_21574, n_21579, n_21580,
       n_21591;
  wire n_21592, n_21593, n_21594, n_21595, n_21598, n_21601, n_21606,
       n_21607;
  wire n_21612, n_21613, n_21618, n_21619, n_21624, n_21625, n_21630,
       n_21631;
  wire n_21636, n_21637, n_21642, n_21643, n_21648, n_21652, n_21657,
       n_21658;
  wire n_21661, n_21664, n_21671, n_21672, n_21673, n_21678, n_21679,
       n_21684;
  wire n_21685, n_21690, n_21691, n_21696, n_21697, n_21702, n_21703,
       n_21708;
  wire n_21709, n_21714, n_21715, n_21720, n_21721, n_21726, n_21727,
       n_21732;
  wire n_21733, n_21744, n_21745, n_21746, n_21747, n_21748, n_21753,
       n_21754;
  wire n_21757, n_21760, n_21765, n_21766, n_21771, n_21772, n_21777,
       n_21778;
  wire n_21783, n_21784, n_21789, n_21790, n_21801, n_21802, n_21803,
       n_21804;
  wire n_21805, n_21808, n_21813, n_21814, n_21817, n_21828, n_21829,
       n_21830;
  wire n_21831, n_21832, n_21837, n_21838, n_21841, n_21846, n_21847,
       n_21852;
  wire n_21853, n_21856, n_21859, n_21862, n_21869, n_21870, n_21871,
       n_21876;
  wire n_21877, n_21882, n_21883, n_21888, n_21889, n_21894, n_21895,
       n_21900;
  wire n_21901, n_21906, n_21907, n_21912, n_21913, n_21918, n_21919,
       n_21924;
  wire n_21925, n_21930, n_21931, n_21936, n_21937, n_21942, n_21943,
       n_21950;
  wire n_21951, n_21952, n_21957, n_21958, n_21961, n_21964, n_21967,
       n_21972;
  wire n_21973, n_21976, n_21981, n_21982, n_21987, n_21988, n_21991,
       n_22002;
  wire n_22003, n_22004, n_22005, n_22006, n_22009, n_22012, n_22017,
       n_22018;
  wire n_22023, n_22024, n_22029, n_22041, n_22042, n_22043, n_22044,
       n_22045;
  wire n_22048, n_22051, n_22054, n_22059, n_22060, n_22065, n_22066,
       n_22071;
  wire n_22072, n_22077, n_22078, n_22085, n_22086, n_22087, n_22090,
       n_22093;
  wire n_22098, n_22099, n_22110, n_22111, n_22112, n_22113, n_22114,
       n_22119;
  wire n_22120, n_22127, n_22128, n_22129, n_22134, n_22135, n_22140,
       n_22141;
  wire n_22146, n_22147, n_22152, n_22153, n_22158, n_22159, n_22164,
       n_22165;
  wire n_22170, n_22171, n_22176, n_22177, n_22184, n_22185, n_22186,
       n_22191;
  wire n_22192, n_22197, n_22198, n_22203, n_22204, n_22209, n_22213,
       n_22216;
  wire n_22219, n_22224, n_22232, n_22233, n_22234, n_22237, n_22240,
       n_22243;
  wire n_22248, n_22249, n_22252, n_22257, n_22258, n_22265, n_22266,
       n_22267;
  wire n_22270, n_22273, n_22278, n_22279, n_22284, n_22285, n_22290,
       n_22291;
  wire n_22296, n_22297, n_22302, n_22303, n_22308, n_22309, n_22314,
       n_22315;
  wire n_22320, n_22321, n_22326, n_22327, n_22332, n_22333, n_22336,
       n_22339;
  wire n_22342, n_22349, n_22350, n_22351, n_22356, n_22357, n_22362,
       n_22363;
  wire n_22368, n_22369, n_22374, n_22375, n_22380, n_22381, n_22386,
       n_22387;
  wire n_22392, n_22393, n_22398, n_22399, n_22406, n_22407, n_22408,
       n_22411;
  wire n_22418, n_22419, n_22420, n_22423, n_22428, n_22429, n_22446,
       n_22447;
  wire n_22448, n_22449, n_22450, n_22451, n_22452, n_22453, n_22456,
       n_22463;
  wire n_22464, n_22465, n_22468, n_22471, n_22478, n_22479, n_22480,
       n_22485;
  wire n_22486, n_22491, n_22492, n_22497, n_22498, n_22503, n_22504,
       n_22509;
  wire n_22510, n_22515, n_22516, n_22521, n_22522, n_22527, n_22528,
       n_22535;
  wire n_22536, n_22537, n_22540, n_22543, n_22546, n_22549, n_22552,
       n_22555;
  wire n_22558, n_22561, n_22564, n_22567, n_22570, n_22573, n_22576,
       n_22579;
  wire n_22582, n_22585, n_22588, n_22591, n_22594, n_22597, n_22600,
       n_22603;
  wire n_22606, n_22609, n_22612, n_22615, n_22618, n_22621, n_22624,
       n_22627;
  wire n_22630, n_22633, n_22638, n_22639, n_22646, n_22647, n_22648,
       n_22656;
  wire n_22657, n_22664, n_22666, n_22669, n_22672, n_22677, n_22678,
       n_22683;
  wire n_22684, n_22689, n_22690, n_22695, n_22696, n_22701, n_22702,
       n_22707;
  wire n_22708, n_22713, n_22714, n_22719, n_22720, n_22725, n_22726,
       n_22731;
  wire n_22732, n_22737, n_22738, n_22743, n_22744, n_22749, n_22750,
       n_22755;
  wire n_22756, n_22761, n_22762, n_22767, n_22768, n_22773, n_22774,
       n_22779;
  wire n_22780, n_22785, n_22786, n_22791, n_22792, n_22797, n_22798,
       n_22803;
  wire n_22804, n_22809, n_22810, n_22815, n_22816, n_22821, n_22822,
       n_22830;
  wire n_22834, n_22837, n_22842, n_22843, n_22848, n_22849, n_22854,
       n_22855;
  wire n_22860, n_22861, n_22866, n_22867, n_22872, n_22873, n_22878,
       n_22879;
  wire n_22884, n_22885, n_22890, n_22891, n_22896, n_22897, n_22902,
       n_22903;
  wire n_22908, n_22909, n_22914, n_22915, n_22920, n_22921, n_22926,
       n_22927;
  wire n_22932, n_22933, n_22938, n_22939, n_22944, n_22945, n_22950,
       n_22951;
  wire n_22956, n_22957, n_22962, n_22963, n_22968, n_22969, n_22974,
       n_22975;
  wire n_22980, n_22981, n_22984, n_22987, n_22990, n_22993, n_22996,
       n_22999;
  wire n_23002, n_23005, n_23008, n_23013, n_23014, n_23021, n_23022,
       n_23023;
  wire n_23032, n_23033, n_23034, n_23035, n_23038, n_23041, n_23044,
       n_23047;
  wire n_23050, n_23053, n_23056, n_23059, n_23062, n_23065, n_23068,
       n_23071;
  wire n_23074, n_23077, n_23080, n_23083, n_23086, n_23089, n_23092,
       n_23095;
  wire n_23098, n_23101, n_23104, n_23107, n_23110, n_23113, n_23116,
       n_23119;
  wire n_23122, n_23125, n_23128, n_23131, n_23134, n_23137, n_23140,
       n_23143;
  wire n_23146, n_23149, n_23152, n_23155, n_23158, n_23161, n_23164,
       n_23167;
  wire n_23170, n_23173, n_23176, n_23179, n_23182, n_23185, n_23188,
       n_23191;
  wire n_23194, n_23197, n_23200, n_23203, n_23206, n_23209, n_23212,
       n_23215;
  wire n_23218, n_23221, n_23224, n_23227, n_23230, n_23233, n_23236,
       n_23239;
  wire n_23242, n_23245, n_23248, n_23251, n_23254, n_23257, n_23260,
       n_23263;
  wire n_23266, n_23269, n_23272, n_23275, n_23278, n_23281, n_23284,
       n_23287;
  wire n_24305, n_24306, n_24307, n_24308, n_24309, n_24310, n_24311,
       n_24312;
  wire n_24313, n_24314, n_24315, n_24316, n_24317, n_24318, n_24319,
       n_24320;
  wire n_24321, n_24322, n_24323, n_24324, n_24325, n_24326, n_24327,
       n_24328;
  wire n_24329, n_24330, n_24331, n_24332, n_24333, n_24334, n_24335,
       n_24336;
  wire n_24339, n_24340, n_24341, n_24342, n_24343, n_24344, n_24345,
       n_24346;
  wire n_24349, n_24350, n_24351, n_24352, n_24353, n_24354, n_24355,
       n_24356;
  wire n_24357, n_24358, n_24359, n_24360, n_24361, n_24362, n_24365,
       n_24366;
  wire n_24367, n_24368, n_24369, n_24370, n_24371, n_24372, n_24373,
       n_24374;
  wire n_24375, n_24376, n_24377, n_24378, n_24379, n_24380, n_24381,
       n_24382;
  wire n_24383, n_24384, n_24385, n_24386, n_24387, n_24388, n_24389,
       n_24390;
  wire n_24391, n_24392, n_24393, n_24394, n_24395, n_24396, n_24397,
       n_24398;
  wire n_24399, n_24400, n_24401, n_24402, n_24403, n_24404, n_24405,
       n_24406;
  wire n_24407, n_24408, n_24411, n_24412, n_24413, n_24414, n_24415,
       n_24416;
  wire n_24417, n_24418, n_24419, n_24420, n_24421, n_24422, n_24423,
       n_24424;
  wire n_24425, n_24426, n_24427, n_24428, n_24429, n_24430, n_24431,
       n_24432;
  wire n_24433, n_24434, n_24435, n_24436, n_24437, n_24438, n_24439,
       n_24440;
  wire n_24441, n_24442, n_24443, n_24444, n_24445, n_24446, n_24447,
       n_24448;
  wire n_24449, n_24450, n_24451, n_24452, n_24453, n_24454, n_24455,
       n_24456;
  wire n_24457, n_24458, n_24459, n_24460, n_24461, n_24462, n_24463,
       n_24464;
  wire n_24465, n_24466, n_24467, n_24468, n_24469, n_24470, n_24471,
       n_24472;
  wire n_24473, n_24474, n_24475, n_24476, n_24477, n_24478, n_24479,
       n_24480;
  wire n_24481, n_24482, n_24483, n_24484, n_24485, n_24486, n_24487,
       n_24488;
  wire n_24489, n_24490, n_24491, n_24492, n_24493, n_24494, n_24495,
       n_24496;
  wire n_24497, n_24498, n_24499, n_24500, n_24501, n_24502, n_24503,
       n_24504;
  wire n_24505, n_24506, n_24507, n_24508, n_24509, n_24510, n_24511,
       n_24512;
  wire n_24513, n_24514, n_24515, n_24516, n_24517, n_24518, n_24519,
       n_24520;
  wire n_24521, n_24523, n_24524, n_24525, n_24526, n_24527, n_24528,
       n_24529;
  wire n_24530, n_24531, n_24532, n_24533, n_24534, n_24535, n_24536,
       n_24537;
  wire n_24538, n_24539, n_24540, n_24541, n_24542, n_24543, n_24544,
       n_24545;
  wire n_24546, n_24547, n_24548, n_24549, n_24550, n_24551, n_24552,
       n_24553;
  wire n_24554, n_24555, n_24556, n_24557, n_24558, n_24559, n_24560,
       n_24561;
  wire n_24562, n_24563, n_24564, n_24565, n_24566, n_24567, n_24568,
       n_24569;
  wire n_24570, n_24571, n_24572, n_24573, n_24574, n_24575, n_24576,
       n_24577;
  wire n_24578, n_24579, n_24580, n_24581, n_24582, n_24583, n_24584,
       n_24585;
  wire n_24586, n_24587, n_24588, n_24589, n_24590, n_24591, n_24592,
       n_24593;
  wire n_24594, n_24595, n_24596, n_24597, n_24598, n_24599, n_24600,
       n_24601;
  wire n_24602, n_24603, n_24604, n_24605, n_24606, n_24607, n_24608,
       n_24609;
  wire n_24610, n_24611, n_24612, n_24613, n_24614, n_24615, n_24616,
       n_24617;
  wire n_24618, n_24619, n_24620, n_24621, n_24622, n_24623, n_24624,
       n_24625;
  wire n_24626, n_24627, n_24628, n_24629, n_24630, n_24631, n_24632,
       n_24633;
  wire n_24634, n_24635, n_24636, n_24637, n_24638, n_24639, n_24640,
       n_24641;
  wire n_24642, n_24643, n_24644, n_24645, n_24646, n_24647, n_24648,
       n_24649;
  wire n_24650, n_24651, n_24652, n_24653, n_24654, n_24655, n_24656,
       n_24657;
  wire n_24658, n_24659, n_24660, n_24661, n_24662, n_24663, n_24664,
       n_24665;
  wire n_24666, n_24667, n_24668, n_24669, n_24670, n_24671, n_24672;
  CDN_flop \data_parity_mem_reg[0] (.clk (clk), .d (n_16947), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[0]));
  CDN_flop \data_parity_mem_reg[1] (.clk (clk), .d (n_16961), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[1]));
  CDN_flop \data_parity_mem_reg[2] (.clk (clk), .d (n_16983), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[2]));
  CDN_flop \data_parity_mem_reg[3] (.clk (clk), .d (n_16972), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[3]));
  CDN_flop \data_parity_mem_reg[4] (.clk (clk), .d (n_17036), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[4]));
  CDN_flop \data_parity_mem_reg[5] (.clk (clk), .d (n_17029), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[5]));
  CDN_flop \data_parity_mem_reg[6] (.clk (clk), .d (n_16992), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[6]));
  CDN_flop \data_parity_mem_reg[7] (.clk (clk), .d (n_17015), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[7]));
  CDN_flop \data_parity_mem_reg[8] (.clk (clk), .d (n_17052), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[8]));
  CDN_flop \data_parity_mem_reg[9] (.clk (clk), .d (n_17007), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_parity_mem[9]));
  CDN_flop \data_stack_mem_reg[0][0] (.clk (clk), .d (n_16932), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [0]));
  CDN_flop \data_stack_mem_reg[0][1] (.clk (clk), .d (n_16937), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [1]));
  CDN_flop \data_stack_mem_reg[0][2] (.clk (clk), .d (n_16936), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [2]));
  CDN_flop \data_stack_mem_reg[0][3] (.clk (clk), .d (n_16935), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [3]));
  CDN_flop \data_stack_mem_reg[0][4] (.clk (clk), .d (n_16934), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [4]));
  CDN_flop \data_stack_mem_reg[0][5] (.clk (clk), .d (n_16933), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [5]));
  CDN_flop \data_stack_mem_reg[0][6] (.clk (clk), .d (n_16931), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [6]));
  CDN_flop \data_stack_mem_reg[0][7] (.clk (clk), .d (n_16938), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[0] [7]));
  CDN_flop \data_stack_mem_reg[1][0] (.clk (clk), .d (n_16959), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [0]));
  CDN_flop \data_stack_mem_reg[1][1] (.clk (clk), .d (n_16955), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [1]));
  CDN_flop \data_stack_mem_reg[1][2] (.clk (clk), .d (n_16954), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [2]));
  CDN_flop \data_stack_mem_reg[1][3] (.clk (clk), .d (n_16956), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [3]));
  CDN_flop \data_stack_mem_reg[1][4] (.clk (clk), .d (n_16957), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [4]));
  CDN_flop \data_stack_mem_reg[1][5] (.clk (clk), .d (n_16953), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [5]));
  CDN_flop \data_stack_mem_reg[1][6] (.clk (clk), .d (n_16958), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [6]));
  CDN_flop \data_stack_mem_reg[1][7] (.clk (clk), .d (n_16960), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[1] [7]));
  CDN_flop \data_stack_mem_reg[2][0] (.clk (clk), .d (n_16976), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [0]));
  CDN_flop \data_stack_mem_reg[2][1] (.clk (clk), .d (n_16977), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [1]));
  CDN_flop \data_stack_mem_reg[2][2] (.clk (clk), .d (n_16975), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [2]));
  CDN_flop \data_stack_mem_reg[2][3] (.clk (clk), .d (n_16980), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [3]));
  CDN_flop \data_stack_mem_reg[2][4] (.clk (clk), .d (n_16981), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [4]));
  CDN_flop \data_stack_mem_reg[2][5] (.clk (clk), .d (n_16979), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [5]));
  CDN_flop \data_stack_mem_reg[2][6] (.clk (clk), .d (n_16978), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [6]));
  CDN_flop \data_stack_mem_reg[2][7] (.clk (clk), .d (n_16982), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[2] [7]));
  CDN_flop \data_stack_mem_reg[3][0] (.clk (clk), .d (n_16970), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [0]));
  CDN_flop \data_stack_mem_reg[3][1] (.clk (clk), .d (n_16965), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [1]));
  CDN_flop \data_stack_mem_reg[3][2] (.clk (clk), .d (n_16971), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [2]));
  CDN_flop \data_stack_mem_reg[3][3] (.clk (clk), .d (n_16964), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [3]));
  CDN_flop \data_stack_mem_reg[3][4] (.clk (clk), .d (n_16969), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [4]));
  CDN_flop \data_stack_mem_reg[3][5] (.clk (clk), .d (n_16968), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [5]));
  CDN_flop \data_stack_mem_reg[3][6] (.clk (clk), .d (n_16967), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [6]));
  CDN_flop \data_stack_mem_reg[3][7] (.clk (clk), .d (n_16966), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[3] [7]));
  CDN_flop \data_stack_mem_reg[4][0] (.clk (clk), .d (n_17037), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [0]));
  CDN_flop \data_stack_mem_reg[4][1] (.clk (clk), .d (n_17040), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [1]));
  CDN_flop \data_stack_mem_reg[4][2] (.clk (clk), .d (n_17038), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [2]));
  CDN_flop \data_stack_mem_reg[4][3] (.clk (clk), .d (n_17039), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [3]));
  CDN_flop \data_stack_mem_reg[4][4] (.clk (clk), .d (n_17041), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [4]));
  CDN_flop \data_stack_mem_reg[4][5] (.clk (clk), .d (n_17033), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [5]));
  CDN_flop \data_stack_mem_reg[4][6] (.clk (clk), .d (n_17034), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [6]));
  CDN_flop \data_stack_mem_reg[4][7] (.clk (clk), .d (n_17035), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[4] [7]));
  CDN_flop \data_stack_mem_reg[5][0] (.clk (clk), .d (n_17022), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [0]));
  CDN_flop \data_stack_mem_reg[5][1] (.clk (clk), .d (n_17023), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [1]));
  CDN_flop \data_stack_mem_reg[5][2] (.clk (clk), .d (n_17024), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [2]));
  CDN_flop \data_stack_mem_reg[5][3] (.clk (clk), .d (n_17025), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [3]));
  CDN_flop \data_stack_mem_reg[5][4] (.clk (clk), .d (n_17030), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [4]));
  CDN_flop \data_stack_mem_reg[5][5] (.clk (clk), .d (n_17026), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [5]));
  CDN_flop \data_stack_mem_reg[5][6] (.clk (clk), .d (n_17027), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [6]));
  CDN_flop \data_stack_mem_reg[5][7] (.clk (clk), .d (n_17028), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[5] [7]));
  CDN_flop \data_stack_mem_reg[6][0] (.clk (clk), .d (n_16993), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [0]));
  CDN_flop \data_stack_mem_reg[6][1] (.clk (clk), .d (n_16994), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [1]));
  CDN_flop \data_stack_mem_reg[6][2] (.clk (clk), .d (n_16991), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [2]));
  CDN_flop \data_stack_mem_reg[6][3] (.clk (clk), .d (n_16990), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [3]));
  CDN_flop \data_stack_mem_reg[6][4] (.clk (clk), .d (n_16989), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [4]));
  CDN_flop \data_stack_mem_reg[6][5] (.clk (clk), .d (n_16988), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [5]));
  CDN_flop \data_stack_mem_reg[6][6] (.clk (clk), .d (n_16995), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [6]));
  CDN_flop \data_stack_mem_reg[6][7] (.clk (clk), .d (n_16996), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[6] [7]));
  CDN_flop \data_stack_mem_reg[7][0] (.clk (clk), .d (n_17012), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [0]));
  CDN_flop \data_stack_mem_reg[7][1] (.clk (clk), .d (n_17018), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [1]));
  CDN_flop \data_stack_mem_reg[7][2] (.clk (clk), .d (n_17011), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [2]));
  CDN_flop \data_stack_mem_reg[7][3] (.clk (clk), .d (n_17017), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [3]));
  CDN_flop \data_stack_mem_reg[7][4] (.clk (clk), .d (n_17016), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [4]));
  CDN_flop \data_stack_mem_reg[7][5] (.clk (clk), .d (n_17014), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [5]));
  CDN_flop \data_stack_mem_reg[7][6] (.clk (clk), .d (n_17019), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [6]));
  CDN_flop \data_stack_mem_reg[7][7] (.clk (clk), .d (n_17013), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[7] [7]));
  CDN_flop \data_stack_mem_reg[8][0] (.clk (clk), .d (n_17045), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [0]));
  CDN_flop \data_stack_mem_reg[8][1] (.clk (clk), .d (n_17051), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [1]));
  CDN_flop \data_stack_mem_reg[8][2] (.clk (clk), .d (n_17044), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [2]));
  CDN_flop \data_stack_mem_reg[8][3] (.clk (clk), .d (n_17046), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [3]));
  CDN_flop \data_stack_mem_reg[8][4] (.clk (clk), .d (n_17047), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [4]));
  CDN_flop \data_stack_mem_reg[8][5] (.clk (clk), .d (n_17048), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [5]));
  CDN_flop \data_stack_mem_reg[8][6] (.clk (clk), .d (n_17049), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [6]));
  CDN_flop \data_stack_mem_reg[8][7] (.clk (clk), .d (n_17050), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[8] [7]));
  CDN_flop \data_stack_mem_reg[9][0] (.clk (clk), .d (n_17004), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[9] [0]));
  CDN_flop \data_stack_mem_reg[9][1] (.clk (clk), .d (n_17000), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[9] [1]));
  CDN_flop \data_stack_mem_reg[9][2] (.clk (clk), .d (n_17006), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[9] [2]));
  CDN_flop \data_stack_mem_reg[9][3] (.clk (clk), .d (n_16999), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[9] [3]));
  CDN_flop \data_stack_mem_reg[9][4] (.clk (clk), .d (n_17003), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[9] [4]));
  CDN_flop \data_stack_mem_reg[9][5] (.clk (clk), .d (n_17001), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[9] [5]));
  CDN_flop \data_stack_mem_reg[9][6] (.clk (clk), .d (n_17005), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[9] [6]));
  CDN_flop \data_stack_mem_reg[9][7] (.clk (clk), .d (n_17002), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\data_stack_mem[9] [7]));
  CDN_flop \data_stack_pointer_reg[0] (.clk (clk), .d (n_16140), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[0]));
  CDN_flop \data_stack_pointer_reg[1] (.clk (clk), .d (n_16925), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[1]));
  CDN_flop \data_stack_pointer_reg[2] (.clk (clk), .d (n_17058), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[2]));
  CDN_flop \data_stack_pointer_reg[3] (.clk (clk), .d (n_17060), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[3]));
  CDN_flop \data_stack_pointer_reg[4] (.clk (clk), .d (n_17061), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (data_stack_pointer[4]));
  CDN_flop dout_valid_reg(.clk (clk), .d (n_16106), .sena (1'b1), .aclr
       (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (dout_valid));
  or g21940 (n_16141, data_stack_pointer[3], data_stack_pointer[1]);
  nand g22329 (n_16357, n_16160, \data_stack_mem[2] [3]);
  nand g22366 (n_16436, n_16160, \data_stack_mem[2] [4]);
  nand g22399 (n_16433, n_16158, \data_stack_mem[3] [4]);
  nand g22511 (n_16587, n_16154, \data_stack_mem[5] [6]);
  nand g22553 (n_16266, n_16154, \data_stack_mem[5] [2]);
  nand g22565 (n_16197, n_16154, \data_stack_mem[5] [1]);
  nand g22577 (n_16155, n_16154, \data_stack_mem[5] [0]);
  nand g22656 (n_16778, n_16158, \data_stack_mem[3] [7]);
  nand g22684 (n_16199, n_16158, \data_stack_mem[3] [1]);
  nand g22703 (n_16352, n_16146, \data_stack_mem[8] [3]);
  nand g22710 (n_16772, n_16146, \data_stack_mem[8] [7]);
  or g26406 (n_16928, wc, data_stack_pointer[3]);
  not gc (wc, data_stack_pointer[1]);
  nand g26464 (n_16172, n_16171, \data_stack_mem[9] [0]);
  or g28043 (n_16152, n_16148, wc0);
  not gc0 (wc0, n_16151);
  or g30819 (n_16926, n_16137, data_stack_pointer[0]);
  nand g30837 (n_16245, n_16166, \data_stack_mem[4] [0]);
  nand g30841 (n_16249, \data_stack_mem[2] [0], n_16164);
  nand g30845 (n_16243, n_16167, \data_stack_mem[5] [0]);
  nand g30852 (n_16241, n_16168, \data_stack_mem[6] [0]);
  nand g30856 (n_16238, n_16170, \data_stack_mem[8] [0]);
  nand g30864 (n_16247, n_16165, \data_stack_mem[3] [0]);
  or g30873 (n_16706, n_16696, n_16705);
  or g30874 (n_16804, n_16706, n_16803);
  or g30878 (n_16711, n_16695, n_16710);
  or g30879 (n_16810, n_16711, n_16809);
  nand g30892 (n_16240, n_16169, \data_stack_mem[7] [0]);
  nand g30921 (n_16264, n_16145, \data_stack_mem[9] [2]);
  nand g30931 (n_16195, n_16145, \data_stack_mem[9] [1]);
  nand g30936 (n_16351, n_16145, \data_stack_mem[9] [3]);
  or g30941 (n_16142, n_16141, data_stack_pointer[0]);
  nand g30951 (n_16429, n_16145, \data_stack_mem[9] [4]);
  nand g30956 (n_16586, n_16145, \data_stack_mem[9] [6]);
  nand g30961 (n_16771, n_16145, \data_stack_mem[9] [7]);
  or g30985 (n_16177, sh_reg_in[4], sh_reg_in[5]);
  nand g31000 (n_16150, data_stack_pointer[1], data_stack_pointer[0]);
  or g31003 (n_16160, wc1, n_16158);
  not gc1 (wc1, n_16150);
  nand g31114 (n_16180, \data_stack_mem[1] [0], \data_stack_mem[0] [0]);
  or g31125 (n_16713, n_16694, n_16712);
  or g31135 (n_16709, n_16708, n_16707);
  or g31297 (n_16702, n_16701, n_16700);
  or g31393 (n_16067, n_16066, sh_reg_out_bit_counter[3]);
  or g31394 (n_16068, n_16067, sh_reg_out_bit_counter[4]);
  or g31407 (n_16065, sh_reg_out_bit_counter[0],
       sh_reg_out_bit_counter[1]);
  or g31408 (n_16066, n_16065, sh_reg_out_bit_counter[2]);
  or g31411 (n_16174, sh_reg_in[1], sh_reg_in[0]);
  nand g31432 (n_16501, n_16158, \data_stack_mem[3] [5]);
  nand g31436 (n_16502, \data_stack_mem[5] [5], n_16154);
  nand g31443 (n_16503, n_16160, \data_stack_mem[2] [5]);
  nand g31447 (n_16504, n_16156, \data_stack_mem[4] [5]);
  nand g31456 (n_16505, n_16148, \data_stack_mem[7] [5]);
  nand g31460 (n_16506, n_16152, \data_stack_mem[6] [5]);
  or g31478 (n_16806, n_16805, n_16709);
  or g31517 (n_16704, n_16697, n_16703);
  or g31711 (n_16835, n_16719, n_16714);
  or g31834 (n_16077, sh_bit_cnt[3], n_16076);
  or g32163 (n_16163, wc2, \data_stack_mem[0] [0]);
  not gc2 (wc2, \data_stack_mem[1] [0]);
  or g32182 (n_16151, n_16150, wc3);
  not gc3 (wc3, data_stack_pointer[2]);
  or g32249 (n_16222, n_16165, wc4);
  not gc4 (wc4, \data_stack_mem[3] [0]);
  or g32276 (n_16220, n_16166, wc5);
  not gc5 (wc5, \data_stack_mem[4] [0]);
  or g32302 (n_16218, n_16167, wc6);
  not gc6 (wc6, \data_stack_mem[5] [0]);
  or g32326 (n_16216, n_16168, wc7);
  not gc7 (wc7, \data_stack_mem[6] [0]);
  or g32335 (n_16232, n_16169, wc8);
  not gc8 (wc8, \data_stack_mem[7] [0]);
  or g32368 (n_16214, n_16170, wc9);
  not gc9 (wc9, \data_stack_mem[8] [0]);
  or g32377 (n_16236, n_16171, wc10);
  not gc10 (wc10, \data_stack_mem[9] [0]);
  or g32520 (n_16826, n_16825, wc11);
  not gc11 (wc11, n_16824);
  or g32583 (n_16837, n_16835, n_16836);
  or g32585 (n_16812, n_16713, n_16811);
  not g38470 (n_16074, rst_n);
  not g38471 (n_16075, enable_n);
  not g38472 (n_16080, n_16079);
  not g38473 (n_16082, n_16081);
  not g38474 (n_16085, n_16084);
  not g38475 (n_16087, n_16086);
  not g38476 (n_16089, n_16088);
  not g38477 (n_16091, n_16090);
  not g38478 (n_16093, n_16092);
  not g38479 (n_16095, n_16094);
  or g38513 (n_16137, data_stack_pointer[4], data_stack_pointer[2]);
  nand g38517 (n_16147, n_16146, \data_stack_mem[8] [0]);
  nand g38520 (n_16149, n_16148, \data_stack_mem[7] [0]);
  or g38521 (n_16148, data_stack_pointer[3], data_stack_pointer[4]);
  nand g38523 (n_16153, n_16152, \data_stack_mem[6] [0]);
  nand g38525 (n_16157, n_16156, \data_stack_mem[4] [0]);
  nand g38527 (n_16159, n_16158, \data_stack_mem[3] [0]);
  or g38528 (n_16158, n_16137, data_stack_pointer[3]);
  nand g38530 (n_16161, n_16160, \data_stack_mem[2] [0]);
  or g38531 (n_16162, n_16158, data_stack_pointer[1]);
  or g38533 (n_16181, wc12, \data_stack_mem[2] [0]);
  not gc12 (wc12, n_16160);
  nand g38543 (n_16196, n_16152, \data_stack_mem[6] [1]);
  nand g38545 (n_16200, n_16160, \data_stack_mem[2] [1]);
  nand g38546 (n_16207, n_16156, \data_stack_mem[4] [1]);
  nand g38547 (n_16210, n_16148, \data_stack_mem[7] [1]);
  nand g38548 (n_16212, n_16146, \data_stack_mem[8] [1]);
  or g38549 (n_16224, wc13, \data_stack_mem[2] [1]);
  not gc13 (wc13, n_16160);
  nand g38552 (n_16265, n_16152, \data_stack_mem[6] [2]);
  nand g38553 (n_16268, n_16158, \data_stack_mem[3] [2]);
  nand g38554 (n_16269, n_16156, \data_stack_mem[4] [2]);
  nand g38556 (n_16271, n_16160, \data_stack_mem[2] [2]);
  nand g38557 (n_16279, n_16148, \data_stack_mem[7] [2]);
  nand g38558 (n_16281, n_16146, \data_stack_mem[8] [2]);
  or g38559 (n_16296, wc14, \data_stack_mem[3] [2]);
  not gc14 (wc14, n_16158);
  nand g38575 (n_16353, n_16148, \data_stack_mem[7] [3]);
  nand g38576 (n_16355, n_16154, \data_stack_mem[5] [3]);
  nand g38577 (n_16356, n_16156, \data_stack_mem[4] [3]);
  nand g38579 (n_16364, n_16158, \data_stack_mem[3] [3]);
  nand g38580 (n_16367, n_16152, \data_stack_mem[6] [3]);
  or g38582 (n_16382, wc15, \data_stack_mem[3] [3]);
  not gc15 (wc15, n_16158);
  nand g38592 (n_16430, n_16154, \data_stack_mem[5] [4]);
  nand g38593 (n_16431, n_16152, \data_stack_mem[6] [4]);
  nand g38595 (n_16434, n_16156, \data_stack_mem[4] [4]);
  nand g38597 (n_16444, n_16148, \data_stack_mem[7] [4]);
  nand g38598 (n_16446, n_16146, \data_stack_mem[8] [4]);
  or g38600 (n_16458, wc16, \data_stack_mem[2] [4]);
  not gc16 (wc16, n_16160);
  nand g38621 (n_16588, n_16152, \data_stack_mem[6] [6]);
  nand g38622 (n_16590, n_16158, \data_stack_mem[3] [6]);
  nand g38623 (n_16591, n_16156, \data_stack_mem[4] [6]);
  nand g38625 (n_16593, n_16160, \data_stack_mem[2] [6]);
  nand g38626 (n_16601, n_16148, \data_stack_mem[7] [6]);
  nand g38627 (n_16603, n_16146, \data_stack_mem[8] [6]);
  or g38629 (n_16616, wc17, \data_stack_mem[2] [6]);
  not gc17 (wc17, n_16160);
  nand g38640 (n_16667, n_16148, \data_stack_mem[7] [7]);
  nand g38641 (n_16676, n_16160, \data_stack_mem[2] [7]);
  or g38642 (n_16677, wc18, \data_stack_mem[2] [7]);
  not gc18 (wc18, n_16160);
  nand g38660 (n_16774, n_16154, \data_stack_mem[5] [7]);
  nand g38661 (n_16775, n_16152, \data_stack_mem[6] [7]);
  nand g38662 (n_16777, n_16156, \data_stack_mem[4] [7]);
  or g39235 (n_17053, sh_bit_cnt[0], enable_n);
  or g39395 (n_17265, wc19, n_16164);
  not gc19 (wc19, \data_stack_mem[2] [0]);
  or g39396 (n_16226, n_17265, n_16225);
  or g39462 (n_17293, n_16813, n_16837);
  or g39476 (n_17298, data_stack_pointer[3], data_stack_pointer[2]);
  or g39488 (n_17303, \data_stack_mem[1] [5], \data_stack_mem[0] [5]);
  nand g39503 (n_17310, n_16145, \data_stack_mem[9] [5]);
  or g39526 (n_17315, \data_stack_mem[8] [4], n_16448);
  or g39529 (n_17316, wc20, n_16474);
  not gc20 (wc20, \data_stack_mem[8] [4]);
  nand g39535 (n_17318, \data_stack_mem[5] [7], n_16723);
  or g39538 (n_17319, \data_stack_mem[2] [6], n_16615);
  or g39541 (n_17320, wc21, n_16636);
  not gc21 (wc21, \data_stack_mem[5] [6]);
  or g39544 (n_17321, wc22, n_16492);
  not gc22 (wc22, \data_stack_mem[9] [4]);
  or g39547 (n_17322, wc23, n_16642);
  not gc23 (wc23, \data_stack_mem[2] [6]);
  or g39550 (n_17323, wc24, n_16490);
  not gc24 (wc24, \data_stack_mem[7] [4]);
  or g39553 (n_17324, wc25, n_16390);
  not gc25 (wc25, \data_stack_mem[9] [3]);
  or g39556 (n_17325, \data_stack_mem[9] [3], n_16414);
  or g39562 (n_17327, wc26, n_16289);
  not gc26 (wc26, \data_stack_mem[4] [2]);
  or g39565 (n_17328, \data_stack_mem[6] [1], wc27);
  not gc27 (wc27, n_16241);
  or g39571 (n_17330, \data_stack_mem[5] [6], n_16609);
  or g39574 (n_17331, wc28, n_16513);
  not gc28 (wc28, \data_stack_mem[5] [5]);
  or g39577 (n_17332, \data_stack_mem[6] [5], n_16547);
  or g39580 (n_17333, wc29, n_16370);
  not gc29 (wc29, \data_stack_mem[8] [3]);
  or g39583 (n_17334, \data_stack_mem[8] [3], n_16394);
  nand g39589 (n_17336, \data_stack_mem[4] [7], n_16725);
  or g39592 (n_17337, wc30, n_16638);
  not gc30 (wc30, \data_stack_mem[4] [6]);
  or g39595 (n_17338, \data_stack_mem[6] [4], n_16450);
  or g39598 (n_17339, \data_stack_mem[5] [5], n_16549);
  or g39601 (n_17340, wc31, n_16476);
  not gc31 (wc31, \data_stack_mem[6] [4]);
  or g39604 (n_17341, wc32, n_16388);
  not gc32 (wc32, \data_stack_mem[7] [3]);
  or g39607 (n_17342, \data_stack_mem[7] [3], n_16412);
  or g39610 (n_17343, \data_stack_mem[9] [2], n_16329);
  or g39613 (n_17344, wc33, n_16305);
  not gc33 (wc33, \data_stack_mem[9] [2]);
  or g39622 (n_17347, wc34, n_16377);
  not gc34 (wc34, \data_stack_mem[2] [3]);
  or g39625 (n_17348, wc35, n_16220);
  not gc35 (wc35, \data_stack_mem[4] [1]);
  or g39631 (n_17350, \data_stack_mem[2] [4], n_16461);
  or g39634 (n_17351, wc36, n_16372);
  not gc36 (wc36, \data_stack_mem[6] [3]);
  or g39637 (n_17352, wc37, n_16515);
  not gc37 (wc37, \data_stack_mem[4] [5]);
  or g39646 (n_17355, \data_stack_mem[6] [3], n_16396);
  or g39652 (n_17357, \data_stack_mem[8] [2], n_16309);
  or g39655 (n_17358, wc38, n_16283);
  not gc38 (wc38, \data_stack_mem[8] [2]);
  or g39661 (n_17360, wc39, n_16678);
  not gc39 (wc39, \data_stack_mem[2] [7]);
  or g39664 (n_17361, \data_stack_mem[7] [6], n_16625);
  nand g39667 (n_17362, \data_stack_mem[3] [7], n_16727);
  or g39670 (n_17363, \data_stack_mem[5] [4], n_16452);
  or g39673 (n_17364, \data_stack_mem[4] [5], n_16551);
  or g39676 (n_17365, wc40, n_16291);
  not gc40 (wc40, \data_stack_mem[2] [2]);
  or g39679 (n_17366, n_16757, n_16758);
  or g39686 (n_17369, \data_stack_mem[1] [1], \data_stack_mem[0] [1]);
  or g39695 (n_17372, wc41, n_16236);
  not gc41 (wc41, \data_stack_mem[9] [1]);
  or g39698 (n_17373, data_stack_pointer[0], n_16928);
  nand g39701 (n_17374, \data_stack_mem[2] [7], n_16729);
  or g39704 (n_17375, wc42, n_16517);
  not gc42 (wc42, \data_stack_mem[3] [5]);
  or g39707 (n_17376, \data_stack_mem[6] [2], n_16311);
  or g39710 (n_17377, \data_stack_mem[3] [6], n_16613);
  or g39713 (n_17378, \data_stack_mem[2] [2], n_16317);
  or g39716 (n_17379, wc43, n_16374);
  not gc43 (wc43, \data_stack_mem[5] [3]);
  or g39719 (n_17380, \data_stack_mem[5] [3], n_16398);
  or g39722 (n_17381, wc44, n_16285);
  not gc44 (wc44, \data_stack_mem[6] [2]);
  or g39728 (n_17383, wc45, n_16287);
  not gc45 (wc45, \data_stack_mem[5] [2]);
  or g39731 (n_17384, \data_stack_mem[2] [1], wc46);
  not gc46 (wc46, n_16249);
  or g39734 (n_17385, wc47, n_16652);
  not gc47 (wc47, \data_stack_mem[9] [6]);
  or g39737 (n_17386, \data_stack_mem[5] [2], n_16313);
  or g39740 (n_17387, wc48, n_16926);
  not gc48 (wc48, data_stack_pointer[3]);
  or g39743 (n_17388, wc49, n_16508);
  not gc49 (wc49, \data_stack_mem[8] [5]);
  or g39746 (n_17389, wc50, n_16532);
  not gc50 (wc50, \data_stack_mem[9] [5]);
  or g39752 (n_17391, \data_stack_mem[1] [3], \data_stack_mem[0] [3]);
  or g39755 (n_17392, n_16826, wc51);
  not gc51 (wc51, n_16829);
  or g39758 (n_17393, wc52, n_16255);
  not gc52 (wc52, n_16240);
  or g39761 (n_17394, wc53, n_16232);
  not gc53 (wc53, \data_stack_mem[7] [1]);
  or g39764 (n_17395, \data_stack_mem[3] [4], n_16456);
  or g39767 (n_17396, \data_stack_mem[8] [6], n_16605);
  or g39770 (n_17397, wc54, n_16216);
  not gc54 (wc54, \data_stack_mem[6] [1]);
  or g39773 (n_17398, wc55, n_16519);
  not gc55 (wc55, \data_stack_mem[2] [5]);
  or g39776 (n_17399, wc56, n_16383);
  not gc56 (wc56, \data_stack_mem[3] [3]);
  or g39779 (n_17400, \data_stack_mem[4] [3], n_16400);
  or g39784 (n_17402, \data_stack_mem[3] [5], n_16553);
  or g39787 (n_17403, \data_stack_mem[2] [5], n_16555);
  or g39790 (n_17404, wc57, n_16484);
  not gc57 (wc57, \data_stack_mem[2] [4]);
  or g39793 (n_17405, wc58, n_16218);
  not gc58 (wc58, \data_stack_mem[5] [1]);
  or g39796 (n_17406, \data_stack_mem[3] [3], n_16407);
  or g39799 (n_17407, \data_stack_mem[4] [2], n_16315);
  or g39802 (n_17408, wc59, n_16297);
  not gc59 (wc59, \data_stack_mem[3] [2]);
  or g39805 (n_17409, \data_stack_mem[5] [1], wc60);
  not gc60 (wc60, n_16243);
  or g39814 (n_17412, wc61, n_16631);
  not gc61 (wc61, \data_stack_mem[8] [6]);
  or g39817 (n_17413, \data_stack_mem[4] [6], n_16611);
  or g39820 (n_17414, \data_stack_mem[3] [2], n_16322);
  or g39823 (n_17415, \data_stack_mem[4] [1], wc62);
  not gc62 (wc62, n_16245);
  or g39829 (n_17417, \data_stack_mem[1] [2], \data_stack_mem[0] [2]);
  or g39832 (n_17418, wc63, n_16640);
  not gc63 (wc63, \data_stack_mem[3] [6]);
  or g39840 (n_17421, wc64, n_16214);
  not gc64 (wc64, \data_stack_mem[8] [1]);
  or g39843 (n_17422, \data_stack_mem[8] [1], wc65);
  not gc65 (wc65, n_16238);
  or g39846 (n_17423, \data_stack_mem[8] [5], n_16543);
  or g39854 (n_17426, n_16649, n_16633);
  or g39857 (n_17427, \data_stack_mem[1] [6], \data_stack_mem[0] [6]);
  or g39862 (n_17429, \data_stack_mem[3] [1], wc66);
  not gc66 (wc66, n_16247);
  or g39868 (n_17431, n_16326, n_16327);
  nand g39879 (n_17435, \data_stack_mem[8] [7], n_16720);
  or g39885 (n_17437, \data_stack_mem[9] [6], n_16629);
  or g39888 (n_17438, wc67, n_16691);
  not gc67 (wc67, \data_stack_mem[7] [7]);
  or g39897 (n_17441, \data_stack_mem[9] [4], n_16470);
  or g39906 (n_17444, \data_stack_mem[2] [3], n_16402);
  or g39909 (n_17445, n_16466, n_16468);
  or g39912 (n_17446, wc68, n_16303);
  not gc68 (wc68, \data_stack_mem[7] [2]);
  or g39915 (n_17447, \data_stack_mem[1] [4], \data_stack_mem[0] [4]);
  or g39921 (n_17449, wc69, n_16634);
  not gc69 (wc69, \data_stack_mem[6] [6]);
  or g39924 (n_17450, wc70, n_16222);
  not gc70 (wc70, \data_stack_mem[3] [1]);
  or g39929 (n_17452, \data_stack_mem[4] [4], n_16454);
  nand g39935 (n_17454, \data_stack_mem[6] [7], n_16721);
  or g39937 (n_16722, wc71, n_17430);
  not gc71 (wc71, n_17454);
  or g39940 (n_17456, n_16566, \data_stack_mem[9] [5]);
  or g39943 (n_17457, wc72, n_16480);
  not gc72 (wc72, \data_stack_mem[3] [4]);
  or g39950 (n_16715, wc73, n_17356);
  not gc73 (wc73, n_17459);
  or g39951 (n_17460, \data_stack_mem[7] [5], n_16545);
  nand g39954 (n_17461, n_16146, \data_stack_mem[8] [5]);
  nand g39957 (n_17462, \data_stack_mem[7] [7], n_16738);
  or g39962 (n_17464, wc74, n_16510);
  not gc74 (wc74, \data_stack_mem[7] [5]);
  or g39967 (n_16671, wc75, n_17317);
  not gc75 (wc75, n_17465);
  or g39968 (n_17466, \data_stack_mem[6] [6], n_16607);
  or g39971 (n_17353, wc76, \data_stack_mem[0] [1]);
  not gc76 (wc76, \data_stack_mem[1] [1]);
  or g39972 (n_17442, wc77, \data_stack_mem[0] [2]);
  not gc77 (wc77, \data_stack_mem[1] [2]);
  or g39973 (n_17411, wc78, \data_stack_mem[0] [3]);
  not gc78 (wc78, \data_stack_mem[1] [3]);
  or g39974 (n_17416, wc79, \data_stack_mem[0] [4]);
  not gc79 (wc79, \data_stack_mem[1] [4]);
  or g39975 (n_17425, wc80, \data_stack_mem[0] [5]);
  not gc80 (wc80, \data_stack_mem[1] [5]);
  or g39976 (n_17443, wc81, \data_stack_mem[0] [6]);
  not gc81 (wc81, \data_stack_mem[1] [6]);
  or g39977 (n_17294, \data_stack_mem[1] [7], wc82);
  not gc82 (wc82, \data_stack_mem[0] [7]);
  or g39988 (n_17290, n_16103, wc83);
  not gc83 (wc83, out_fifo_read_pointer[1]);
  or g39989 (n_17300, n_16103, wc84);
  not gc84 (wc84, out_fifo_read_pointer[0]);
  or g40120 (n_17370, wc85, \data_stack_mem[9] [1]);
  not gc85 (wc85, n_16172);
  or g40216 (n_17349, n_16674, wc86);
  not gc86 (wc86, \data_stack_mem[3] [7]);
  or g40226 (n_16728, n_17448, wc87);
  not gc87 (wc87, n_17362);
  or g40238 (n_17329, n_16672, wc88);
  not gc88 (wc88, \data_stack_mem[4] [7]);
  or g40240 (n_16818, n_16746, wc89);
  not gc89 (wc89, n_16749);
  or g40251 (n_16726, n_17345, wc90);
  not gc90 (wc90, n_17336);
  or g40259 (n_17465, n_16670, wc91);
  not gc91 (wc91, \data_stack_mem[5] [7]);
  or g40271 (n_16724, n_17326, wc92);
  not gc92 (wc92, n_17318);
  or g40278 (n_17433, n_16668, wc93);
  not gc93 (wc93, \data_stack_mem[6] [7]);
  or g40295 (n_17459, n_16666, wc94);
  not gc94 (wc94, \data_stack_mem[8] [7]);
  or g40309 (n_17432, n_16717, wc95);
  not gc95 (wc95, \data_stack_mem[9] [7]);
  or g40310 (n_16756, n_17436, wc96);
  not gc96 (wc96, n_17435);
  or g40313 (n_17440, n_16814, wc97);
  not gc97 (wc97, n_16823);
  or g40326 (n_16832, n_16760, wc98);
  not gc98 (wc98, n_16831);
  nand g40479 (n_17481, n_16757, n_16758);
  or g40533 (n_17507, wc99, n_16376);
  not gc99 (wc99, \data_stack_mem[4] [3]);
  or g40536 (n_17508, wc100, n_16478);
  not gc100 (wc100, \data_stack_mem[5] [4]);
  or g40541 (n_17510, wc101, n_16479);
  not gc101 (wc101, \data_stack_mem[4] [4]);
  or g40581 (n_16819, n_16747, wc102);
  not gc102 (wc102, n_16748);
  or g40583 (n_17501, n_16512, wc103);
  not gc103 (wc103, \data_stack_mem[6] [5]);
  nand g40841 (n_17634, \data_stack_mem[9] [7], n_17366);
  nand g40843 (n_17635, \data_stack_mem[1] [0], n_16162);
  or g41013 (n_17720, data_stack_pointer[1], data_stack_pointer[2]);
  nand g41023 (n_17725, \data_stack_mem[9] [0], n_16145);
  or g41041 (n_17734, \data_stack_mem[3] [6], wc104);
  not gc104 (wc104, n_16158);
  or g41045 (n_17736, \data_stack_mem[3] [1], wc105);
  not gc105 (wc105, n_16158);
  nand g41053 (n_17740, n_16162, n_17427);
  nand g41055 (n_17741, n_16162, n_17369);
  or g41057 (n_17742, \data_stack_mem[2] [2], wc106);
  not gc106 (wc106, n_16160);
  or g41061 (n_17744, \data_stack_mem[3] [4], wc107);
  not gc107 (wc107, n_16158);
  or g41065 (n_17746, \data_stack_mem[3] [7], wc108);
  not gc108 (wc108, n_16158);
  nand g41079 (n_17753, n_16162, n_17447);
  nand g41081 (n_17754, n_16162, n_17417);
  or g41083 (n_17755, \data_stack_mem[3] [0], wc109);
  not gc109 (wc109, n_16158);
  or g41089 (n_17758, \data_stack_mem[2] [3], wc110);
  not gc110 (wc110, n_16160);
  nand g41097 (n_17762, n_16162, n_17391);
  or g41121 (n_17716, n_17799, n_17800);
  or g45313 (n_16675, n_17359, wc111);
  not gc111 (wc111, n_17349);
  or g45320 (n_16673, n_17335, wc112);
  not gc112 (wc112, n_17329);
  or g45332 (n_16669, n_17453, wc113);
  not gc113 (wc113, n_17433);
  nand g45356 (n_16890, n_22938, n_22939);
  nand g45357 (n_16891, n_22944, n_22945);
  nand g45358 (n_16892, n_22950, n_22951);
  nand g45359 (n_16897, n_22980, n_22981);
  nand g45360 (n_16894, n_22962, n_22963);
  nand g45361 (n_16895, n_22968, n_22969);
  nand g45362 (n_16896, n_22974, n_22975);
  nand g45363 (n_16893, n_22956, n_22957);
  nand g45372 (n_16857, n_22902, n_22903);
  nand g45373 (n_16855, n_22896, n_22897);
  nand g45374 (n_16861, n_22914, n_22915);
  nand g45375 (n_16863, n_22920, n_22921);
  nand g45376 (n_16853, n_22890, n_22891);
  nand g45377 (n_16865, n_22926, n_22927);
  nand g45378 (n_16867, n_22932, n_22933);
  or g45379 (n_24305, wc114, n_17511);
  not gc114 (wc114, n_17512);
  or g45380 (n_24306, n_17512, wc115);
  not gc115 (wc115, n_17511);
  nand g45381 (n_16889, n_24305, n_24306);
  nand g45382 (n_16859, n_22908, n_22909);
  nand g45383 (n_16842, n_22860, n_22861);
  nand g45384 (n_16876, n_22785, n_22786);
  nand g45385 (n_16843, n_22866, n_22867);
  nand g45386 (n_16877, n_22791, n_22792);
  nand g45387 (n_16875, n_22779, n_22780);
  nand g45388 (n_16844, n_22872, n_22873);
  or g45389 (n_24307, wc116, n_16838);
  not gc116 (wc116, n_16852);
  or g45390 (n_24308, n_16852, wc117);
  not gc117 (wc117, n_16838);
  nand g45391 (n_17512, n_24307, n_24308);
  nand g45392 (n_16845, n_22878, n_22879);
  nand g45393 (n_16841, n_22854, n_22855);
  nand g45394 (n_16846, n_22884, n_22885);
  nand g45395 (n_16878, n_22797, n_22798);
  or g45396 (n_22890, n_16110, n_16852);
  or g45397 (n_22932, n_16131, n_16852);
  nand g45398 (n_16840, n_22848, n_22849);
  nand g45399 (n_16879, n_22803, n_22804);
  or g45400 (n_22926, n_16128, n_16852);
  nand g45401 (n_16839, n_22842, n_22843);
  or g45402 (n_22896, n_16113, n_16852);
  or g45403 (n_22920, n_16125, n_16852);
  nand g45404 (n_16880, n_22809, n_22810);
  nand g45405 (n_16882, n_22821, n_22822);
  or g45406 (n_22914, n_16122, n_16852);
  nand g45407 (n_16881, n_22815, n_22816);
  or g45408 (n_22902, n_16852, n_16116);
  or g45409 (n_22908, n_16119, n_16852);
  or g45412 (n_22848, n_16113, n_16838);
  nand g45413 (n_16864, n_22761, n_22762);
  nand g45414 (n_16849, n_22725, n_22726);
  or g45415 (n_22842, n_16110, n_16838);
  nand g45417 (n_16858, n_22743, n_22744);
  or g45419 (n_22884, n_16131, n_16838);
  nand g45420 (n_16862, n_22755, n_22756);
  or g45422 (n_22878, n_16128, n_16838);
  or g45425 (n_22872, n_16125, n_16838);
  nand g45426 (n_16854, n_22731, n_22732);
  or g45428 (n_22866, n_16122, n_16838);
  nand g45429 (n_16866, n_22767, n_22768);
  nand g45430 (n_16860, n_22749, n_22750);
  or g45431 (n_22860, n_16119, n_16838);
  or g45433 (n_22854, n_16838, n_16116);
  nand g45434 (n_16856, n_22737, n_22738);
  nand g45435 (n_17108, n_17107, n_22600);
  nand g45436 (n_17109, n_17107, n_22603);
  nand g45437 (n_17094, n_17092, n_22567);
  nand g45438 (n_17110, n_17107, n_22606);
  nand g45439 (n_17111, n_17107, n_22609);
  nand g45440 (n_17113, n_17112, n_22612);
  nand g45441 (n_17095, n_17092, n_22570);
  nand g45442 (n_17114, n_17112, n_22615);
  nand g45443 (n_17093, n_17092, n_22564);
  nand g45444 (n_17096, n_17092, n_22573);
  nand g45445 (n_17115, n_17112, n_22618);
  nand g45446 (n_17106, n_17102, n_22597);
  nand g45447 (n_17116, n_17112, n_22621);
  nand g45448 (n_17118, n_17117, n_22624);
  nand g45449 (n_17091, n_17087, n_22561);
  nand g45450 (n_17105, n_17102, n_22594);
  nand g45451 (n_17119, n_17117, n_22627);
  nand g45452 (n_17120, n_17117, n_22630);
  nand g45453 (n_17090, n_17087, n_22558);
  or g45454 (n_24309, wc118, n_16848);
  not gc118 (wc118, n_16762);
  or g45455 (n_24310, n_16762, wc119);
  not gc119 (wc119, n_16848);
  nand g45456 (n_17511, n_24309, n_24310);
  nand g45457 (n_17104, n_17102, n_22591);
  nand g45458 (n_17121, n_17117, n_22633);
  nand g45459 (n_17089, n_17087, n_22555);
  nand g45460 (n_17103, n_17102, n_22588);
  nand g45461 (n_16763, n_22677, n_22678);
  nand g45462 (n_16764, n_22683, n_22684);
  nand g45463 (n_17088, n_17087, n_22552);
  nand g45464 (n_16765, n_22689, n_22690);
  nand g45465 (n_17101, n_17097, n_22585);
  nand g45466 (n_16766, n_22695, n_22696);
  nand g45467 (n_16767, n_22701, n_22702);
  nand g45468 (n_17100, n_17097, n_22582);
  nand g45469 (n_22834, n_17636, n_16851);
  nand g45470 (n_17083, n_17082, n_22540);
  nand g45471 (n_16768, n_22707, n_22708);
  or g45472 (n_24311, wc120, n_16873);
  not gc120 (wc120, n_16870);
  or g45473 (n_24312, n_16870, wc121);
  not gc121 (wc121, n_16873);
  nand g45474 (n_16874, n_24311, n_24312);
  nand g45475 (n_17086, n_17082, n_22549);
  nand g45476 (n_17098, n_17097, n_22576);
  nand g45477 (n_16769, n_22713, n_22714);
  nand g45478 (n_17099, n_17097, n_22579);
  nand g45479 (n_16770, n_22719, n_22720);
  or g45480 (n_22767, n_16131, n_16848);
  or g45481 (n_22725, n_16110, n_16848);
  or g45482 (n_22761, n_16128, n_16848);
  nand g45483 (n_17085, n_17082, n_22546);
  or g45484 (n_22755, n_16125, n_16848);
  or g45485 (n_22731, n_16113, n_16848);
  or g45486 (n_22749, n_16122, n_16848);
  nand g45487 (n_17084, n_17082, n_22543);
  or g45488 (n_22743, n_16119, n_16848);
  or g45489 (n_22737, n_16848, n_16116);
  nand g45491 (n_22837, n_17643, n_16834);
  nand g45492 (n_16793, n_22491, n_22492);
  or g45493 (n_17092, n_17081, n_16090);
  nand g45494 (n_16797, n_22515, n_22516);
  nand g45495 (n_16792, n_22485, n_22486);
  or g45496 (n_22719, n_16131, n_16762);
  nand g45498 (n_24313, n_16868, n_16869);
  or g45499 (n_24314, n_16868, n_16869);
  nand g45500 (n_16870, n_24313, n_24314);
  or g45501 (n_22713, n_16128, n_16762);
  or g45502 (n_17097, n_17081, n_16094);
  nand g45503 (n_16799, n_22527, n_22528);
  or g45504 (n_22707, n_16125, n_16762);
  nand g45505 (n_16794, n_22497, n_22498);
  or g45506 (n_17117, n_17081, n_16086);
  or g45507 (n_22701, n_16122, n_16762);
  nand g45508 (n_16795, n_22503, n_22504);
  or g45509 (n_17112, n_17081, n_16081);
  or g45510 (n_22695, n_16119, n_16762);
  or g45511 (n_17087, n_17081, n_16092);
  or g45512 (n_22689, n_16762, n_16116);
  nand g45513 (n_16796, n_22509, n_22510);
  or g45514 (n_17107, n_17081, n_16084);
  or g45515 (n_17102, n_17081, n_16088);
  or g45516 (n_22683, n_16113, n_16762);
  or g45517 (n_17636, n_22666, n_16175);
  or g45518 (n_17082, n_17081, n_16079);
  or g45519 (n_22677, n_16110, n_16762);
  nand g45520 (n_16798, n_22521, n_22522);
  or g45521 (n_16834, n_22774, n_16176);
  or g45522 (n_22497, n_16791, n_16116);
  or g45523 (n_17643, n_22648, n_16175);
  or g45524 (n_22521, n_16128, n_16791);
  or g45525 (n_17081, n_16883, wc122);
  not gc122 (wc122, rst_n);
  or g45526 (n_22485, n_16110, n_16791);
  or g45527 (n_22515, n_16125, n_16791);
  or g45528 (n_22503, n_16119, n_16791);
  or g45529 (n_16851, wc123, n_16176);
  not gc123 (wc123, n_22830);
  or g45530 (n_22527, n_16131, n_16791);
  nand g45531 (n_22666, n_22664, n_22428);
  or g45532 (n_22491, n_16113, n_16791);
  or g45533 (n_24315, wc124, n_16791);
  not gc124 (wc124, n_16186);
  or g45534 (n_24316, n_16186, wc125);
  not gc125 (wc125, n_16791);
  nand g45535 (n_16869, n_24315, n_24316);
  or g45536 (n_22509, n_16122, n_16791);
  nand g45537 (n_22669, n_17655, n_16847);
  nand g45539 (n_22672, n_17660, n_16761);
  nand g45540 (n_22648, n_22646, n_22647);
  or g45541 (n_16883, n_22429, n_16175);
  nand g45542 (n_22830, n_16833, n_17392);
  or g45543 (n_22664, n_17293, wc126);
  not gc126 (wc126, n_16850);
  or g45544 (n_17655, n_22657, n_16176);
  or g45545 (n_16847, n_22537, n_16175);
  nand g45547 (n_22774, n_16833, n_22773);
  or g45548 (n_16761, n_22639, n_16176);
  or g45551 (n_22647, wc127, n_16813);
  not gc127 (wc127, n_16837);
  or g45552 (n_22646, n_16837, wc128);
  not gc128 (wc128, n_16813);
  nand g45553 (n_22537, n_22535, n_22536);
  or g45554 (n_22480, n_22478, n_22479);
  or g45555 (n_17660, n_22465, n_16175);
  nand g45556 (n_22657, n_16832, n_22656);
  nand g45558 (n_22465, n_22463, n_22464);
  nand g45559 (n_22639, n_16760, n_22638);
  or g45560 (n_22479, wc129, n_16789);
  not gc129 (wc129, n_16786);
  or g45561 (n_22535, n_16835, wc130);
  not gc130 (wc130, n_16836);
  or g45562 (n_22536, wc131, n_16836);
  not gc131 (wc131, n_16835);
  or g45563 (n_24317, wc132, n_16420);
  not gc132 (wc132, n_16872);
  or g45564 (n_24318, n_16872, wc133);
  not gc133 (wc133, n_16420);
  nand g45565 (n_16873, n_24317, n_24318);
  nand g45566 (n_22478, n_17646, n_16790);
  or g45567 (n_22656, n_16831, wc134);
  not gc134 (wc134, n_16760);
  or g45568 (n_24319, wc135, n_16570);
  not gc135 (wc135, n_16871);
  or g45569 (n_24320, n_16871, wc136);
  not gc136 (wc136, n_16570);
  nand g45570 (n_16872, n_24319, n_24320);
  nand g45571 (n_16658, n_22356, n_22357);
  or g45572 (n_16790, n_22408, n_16175);
  nand g45573 (n_16659, n_22362, n_22363);
  nand g45574 (n_16660, n_22368, n_22369);
  nand g45575 (n_16661, n_22374, n_22375);
  or g45576 (n_16786, n_22453, n_16176);
  nand g45578 (n_16662, n_22380, n_22381);
  nand g45581 (n_16663, n_22386, n_22387);
  nand g45583 (n_16664, n_22392, n_22393);
  nand g45584 (n_16665, n_22398, n_22399);
  nand g45585 (n_22408, n_22406, n_22407);
  or g45586 (n_22453, n_22451, n_22452);
  or g45587 (n_22392, n_16128, n_16657);
  or g45588 (n_24321, wc137, n_16657);
  not gc137 (wc137, n_16262);
  or g45589 (n_24322, n_16262, wc138);
  not gc138 (wc138, n_16657);
  nand g45590 (n_16871, n_24321, n_24322);
  or g45593 (n_22386, n_16125, n_16657);
  or g45594 (n_22362, n_16113, n_16657);
  nand g45595 (n_17439, n_16145, n_22471);
  or g45596 (n_22380, n_16122, n_16657);
  nand g45599 (n_16813, n_24323, n_24324);
  or g45600 (n_22356, n_16110, n_16657);
  or g45601 (n_22374, n_16119, n_16657);
  nand g45602 (n_16836, n_16812, n_22468);
  or g45603 (n_22398, n_16131, n_16657);
  or g45604 (n_22368, n_16657, n_16116);
  nand g45605 (n_22471, n_17634, n_17481);
  nand g45607 (n_16577, n_22308, n_22309);
  nand g45608 (n_22452, n_22449, n_22450);
  nand g45609 (n_22423, n_16716, n_17432);
  nand g45610 (n_16583, n_22326, n_22327);
  nand g45611 (n_16714, n_16713, n_22456);
  nand g45613 (n_22468, n_16713, n_16811);
  nand g45614 (n_16585, n_22332, n_22333);
  nand g45615 (n_16579, n_22314, n_22315);
  nand g45616 (n_16571, n_22290, n_22291);
  nand g45617 (n_22451, n_22447, n_22448);
  nand g45618 (n_16573, n_22296, n_22297);
  or g45619 (n_22406, n_16716, n_17662);
  nand g45620 (n_16575, n_22302, n_22303);
  nand g45621 (n_16581, n_22320, n_22321);
  nand g45622 (n_22407, n_17662, n_16716);
  nand g45623 (n_24325, n_16826, n_16829);
  or g45624 (n_24326, n_16826, n_16829);
  nand g45625 (n_16830, n_24325, n_24326);
  nand g45626 (n_22456, n_16712, n_16694);
  or g45628 (n_22290, n_16110, n_16570);
  or g45629 (n_22296, n_16113, n_16570);
  or g45630 (n_22302, n_16570, n_16116);
  or g45631 (n_22308, n_16119, n_16570);
  or g45632 (n_22332, n_16131, n_16570);
  or g45633 (n_22314, n_16122, n_16570);
  or g45634 (n_22450, n_22446, n_16758);
  or g45635 (n_22320, n_16125, n_16570);
  or g45636 (n_22326, n_16128, n_16570);
  or g45637 (n_22449, n_16785, n_17481);
  or g45638 (n_22448, \data_stack_mem[9] [7], n_17366);
  nand g45639 (n_24327, n_16715, n_16693);
  or g45640 (n_24328, n_16715, n_16693);
  nand g45641 (n_16716, n_24327, n_24328);
  or g45642 (n_22351, n_22349, n_22350);
  or g45643 (n_16694, n_17356, wc139);
  not gc139 (wc139, n_22342);
  nand g45646 (n_17284, n_24329, n_24330);
  nand g45647 (n_16811, n_16810, n_22411);
  or g45649 (n_22350, wc140, n_16656);
  not gc140 (wc140, n_16630);
  nand g45650 (n_24331, n_16825, n_16824);
  or g45651 (n_24332, n_16825, n_16824);
  nand g45652 (n_16831, n_24331, n_24332);
  nand g45653 (n_22349, n_17668, n_16653);
  or g45654 (n_22447, n_16757, wc141);
  not gc141 (wc141, n_17645);
  nand g45655 (n_16718, n_16145, n_22270);
  nand g45657 (n_17662, n_22257, n_22258);
  or g45658 (n_16630, n_22267, n_16176);
  nand g45659 (n_22411, n_16711, n_16809);
  nand g45660 (n_24333, n_16756, n_16740);
  or g45661 (n_24334, n_16756, n_16740);
  nand g45662 (n_16757, n_24333, n_24334);
  nand g45663 (n_17356, n_16146, n_22240);
  or g45664 (n_16653, n_22234, n_16175);
  or g45665 (n_22285, wc142, n_22284);
  not gc142 (wc142, n_17424);
  nand g45666 (n_24335, n_16741, n_16754);
  or g45667 (n_24336, n_16741, n_16754);
  nand g45668 (n_16755, n_24335, n_24336);
  nand g45669 (n_17645, n_16145, n_22336);
  nand g45670 (n_16712, n_16711, n_22339);
  or g45671 (n_22270, \data_stack_mem[9] [7], wc143);
  not gc143 (wc143, n_16717);
  or g45672 (n_22257, n_16785, n_16717);
  or g45673 (n_22258, n_16771, wc144);
  not gc144 (wc144, n_16717);
  nand g45674 (n_22342, n_17459, n_16693);
  nand g45675 (n_22267, n_22265, n_22266);
  nand g45676 (n_16717, n_22209, n_23284);
  nand g45677 (n_22339, n_16710, n_16695);
  or g45678 (n_16741, n_17436, wc145);
  not gc145 (wc145, n_22273);
  nand g45679 (n_16693, n_22278, n_22279);
  nand g45680 (n_16584, n_22176, n_22177);
  nand g45684 (n_22234, n_22232, n_22233);
  nand g45685 (n_16582, n_22170, n_22171);
  nand g45686 (n_16580, n_22164, n_22165);
  nand g45688 (n_16499, n_22134, n_22135);
  nand g45689 (n_16578, n_22158, n_22159);
  nand g45690 (n_16572, n_22140, n_22141);
  nand g45691 (n_22336, \data_stack_mem[9] [7], n_16758);
  nand g45692 (n_16576, n_22152, n_22153);
  nand g45693 (n_16574, n_22146, n_22147);
  or g45694 (n_22240, \data_stack_mem[8] [7], wc146);
  not gc146 (wc146, n_16666);
  or g45695 (n_22146, n_16498, n_16116);
  or g45696 (n_22152, n_16119, n_16498);
  or g45697 (n_22158, n_16122, n_16498);
  or g45699 (n_22140, n_16113, n_16498);
  nand g45702 (n_16808, n_24339, n_24340);
  or g45703 (n_22134, n_16110, n_16498);
  or g45705 (n_22164, n_16125, n_16498);
  or g45706 (n_22170, n_16128, n_16498);
  nand g45707 (n_22233, n_17678, n_16651);
  nand g45708 (n_24341, n_16814, n_16823);
  or g45709 (n_24342, n_16814, n_16823);
  nand g45710 (n_16824, n_24341, n_24342);
  or g45711 (n_22232, n_16651, n_17678);
  or g45712 (n_22176, n_16131, n_16498);
  or g45713 (n_22265, n_16627, n_17667);
  nand g45714 (n_22266, n_17667, n_16627);
  nand g45715 (n_24343, n_16335, n_16498);
  or g45716 (n_24344, n_16335, n_16498);
  nand g45717 (n_16868, n_24343, n_24344);
  nand g45718 (n_23284, n_16651, n_17385);
  nand g45720 (n_17436, n_16146, n_22243);
  nand g45721 (n_16758, n_22224, n_23287);
  or g45722 (n_22273, wc147, n_16740);
  not gc147 (wc147, n_17435);
  nand g45723 (n_16569, n_17689, n_16568);
  nand g45724 (n_16666, n_22065, n_23278);
  or g45725 (n_16568, n_22186, n_16176);
  nand g45727 (n_16740, n_22248, n_22249);
  or g45728 (n_22243, \data_stack_mem[8] [7], n_16720);
  nand g45729 (n_24345, n_16742, n_16753);
  or g45730 (n_24346, n_16742, n_16753);
  nand g45731 (n_16754, n_24345, n_24346);
  nand g45732 (n_23287, n_16627, n_17437);
  nand g45733 (n_22252, n_16689, n_17438);
  nand g45734 (n_17667, n_22203, n_22204);
  nand g45735 (n_16809, n_16806, n_22237);
  nand g45739 (n_16692, n_16148, n_22213);
  nand g45740 (n_24349, n_16632, n_16650);
  or g45741 (n_24350, n_16632, n_16650);
  nand g45742 (n_16651, n_24349, n_24350);
  nand g45745 (n_16807, n_24351, n_24352);
  nand g45746 (n_17658, n_22197, n_22198);
  nand g45747 (n_23278, n_17412, n_16650);
  or g45749 (n_22213, \data_stack_mem[7] [7], wc148);
  not gc148 (wc148, n_16691);
  or g45750 (n_22129, n_22127, n_22128);
  or g45751 (n_16742, n_16739, wc149);
  not gc149 (wc149, n_22219);
  nand g45752 (n_24353, n_16606, n_16626);
  or g45753 (n_24354, n_16606, n_16626);
  nand g45754 (n_16627, n_24353, n_24354);
  nand g45755 (n_22224, \data_stack_mem[9] [6], n_16629);
  or g45756 (n_22203, n_16586, n_16629);
  or g45758 (n_22198, n_16667, wc150);
  not gc150 (wc150, n_16691);
  nand g45759 (n_16720, n_22191, n_23281);
  nand g45760 (n_17678, n_22077, n_22078);
  nand g45761 (n_22186, n_22184, n_22185);
  nand g45762 (n_22237, n_16709, n_16805);
  nand g45763 (n_16710, n_16709, n_22216);
  or g45764 (n_16650, wc151, n_22114);
  not gc151 (wc151, n_22113);
  or g45765 (n_17690, n_22087, n_16175);
  nand g45766 (n_24355, n_16815, n_16822);
  or g45767 (n_24356, n_16815, n_16822);
  nand g45768 (n_16823, n_24355, n_24356);
  or g45769 (n_22197, n_16690, n_16691);
  nand g45772 (n_24357, n_16669, n_16688);
  or g45773 (n_24358, n_16669, n_16688);
  nand g45774 (n_16689, n_24357, n_24358);
  nand g45775 (n_22113, n_17651, n_16649);
  or g45777 (n_16632, n_22066, wc152);
  not gc152 (wc152, n_16146);
  or g45778 (n_22077, n_16628, n_16652);
  or g45779 (n_22078, n_16586, wc153);
  not gc153 (wc153, n_16652);
  nand g45780 (n_22216, n_16707, n_16708);
  nand g45781 (n_23281, n_17396, n_16626);
  or g45782 (n_22128, wc154, n_16497);
  not gc154 (wc154, n_16473);
  nand g45783 (n_24359, n_16743, n_16752);
  or g45784 (n_24360, n_16743, n_16752);
  nand g45785 (n_16753, n_24359, n_24360);
  or g45786 (n_22209, \data_stack_mem[9] [6], wc155);
  not gc155 (wc155, n_16652);
  nand g45787 (n_16629, n_22059, n_23275);
  nand g45789 (n_16691, n_22119, n_22120);
  nand g45790 (n_16739, n_16148, n_22090);
  nand g45791 (n_17647, n_22071, n_22072);
  nand g45792 (n_22087, n_22085, n_22086);
  or g45793 (n_16606, n_22192, wc156);
  not gc156 (wc156, n_16146);
  nand g45794 (n_22114, n_22111, n_22112);
  or g45796 (n_22071, n_16667, n_16738);
  or g45797 (n_22119, \data_stack_mem[7] [6], wc157);
  not gc157 (wc157, n_17426);
  nand g45798 (n_24361, n_16722, n_16736);
  or g45799 (n_24362, n_16722, n_16736);
  nand g45800 (n_16737, n_24361, n_24362);
  or g45801 (n_22090, \data_stack_mem[7] [7], n_16738);
  or g45802 (n_16743, n_17430, wc158);
  not gc158 (wc158, n_22051);
  or g45803 (n_16473, n_22045, n_16176);
  nand g45804 (n_16805, n_16804, n_22093);
  nand g45805 (n_22127, n_17695, n_16494);
  or g45806 (n_16567, n_22060, wc159);
  not gc159 (wc159, n_16145);
  or g45807 (n_22112, n_22110, wc160);
  not gc160 (wc160, n_16633);
  or g45808 (n_22111, n_16624, n_17426);
  nand g45812 (n_16827, n_17287, n_17371);
  nand g45813 (n_22066, n_17412, n_22065);
  nand g45815 (n_16652, n_22023, n_23269);
  nand g45816 (n_23275, n_16565, n_17456);
  nand g45817 (n_16626, n_22098, n_22099);
  nand g45820 (n_22192, n_17396, n_22191);
  or g45821 (n_16533, n_22024, wc161);
  not gc161 (wc161, n_16145);
  nand g45822 (n_22054, n_16688, n_17433);
  nand g45823 (n_16707, n_16706, n_22048);
  nand g45824 (n_22060, n_17456, n_22059);
  nand g45825 (n_22120, n_16649, n_16633);
  nand g45826 (n_16738, n_22029, n_23272);
  nand g45829 (n_22093, n_16706, n_16803);
  or g45830 (n_16494, n_22006, n_16175);
  nand g45831 (n_17453, n_16152, n_22009);
  nand g45832 (n_16428, n_21918, n_21919);
  nand g45833 (n_16427, n_21912, n_21913);
  nand g45834 (n_16426, n_21906, n_21907);
  or g45835 (n_22110, n_16649, n_16601);
  nand g45836 (n_24365, n_16816, n_16821);
  or g45837 (n_24366, n_16816, n_16821);
  nand g45838 (n_16822, n_24365, n_24366);
  nand g45839 (n_16425, n_21900, n_21901);
  nand g45840 (n_16424, n_21894, n_21895);
  nand g45841 (n_21952, n_21950, n_21951);
  nand g45842 (n_16423, n_21888, n_21889);
  or g45843 (n_22065, \data_stack_mem[8] [6], wc162);
  not gc162 (wc162, n_16631);
  nand g45844 (n_16422, n_21882, n_21883);
  nand g45845 (n_24367, n_16544, n_16564);
  or g45846 (n_24368, n_16544, n_16564);
  nand g45847 (n_16565, n_24367, n_24368);
  nand g45850 (n_16421, n_21876, n_21877);
  nand g45851 (n_23269, n_16531, n_17389);
  nand g45852 (n_22191, \data_stack_mem[8] [6], n_16605);
  or g45853 (n_21912, n_16128, n_16420);
  or g45854 (n_21882, n_16113, n_16420);
  nand g45855 (n_22048, n_16705, n_16696);
  nand g45856 (n_17430, n_16152, n_22012);
  nand g45857 (n_24369, n_16724, n_16735);
  or g45858 (n_24370, n_16724, n_16735);
  nand g45859 (n_16736, n_24369, n_24370);
  nand g45860 (n_22024, n_17389, n_22023);
  nand g45861 (n_22059, \data_stack_mem[9] [5], n_16566);
  nand g45862 (n_23272, n_16623, n_17361);
  nand g45863 (n_17638, n_21987, n_21988);
  or g45864 (n_21918, n_16131, n_16420);
  nand g45865 (n_24371, n_16509, n_16530);
  or g45866 (n_24372, n_16509, n_16530);
  nand g45867 (n_16531, n_24371, n_24372);
  nand g45868 (n_24373, n_16635, n_16648);
  or g45869 (n_24374, n_16635, n_16648);
  nand g45870 (n_16649, n_24373, n_24374);
  or g45871 (n_21888, n_16420, n_16116);
  or g45872 (n_21894, n_16119, n_16420);
  nand g45873 (n_24375, n_16744, n_16751);
  or g45874 (n_24376, n_16744, n_16751);
  nand g45875 (n_16752, n_24375, n_24376);
  nand g45876 (n_22044, n_22041, n_22042);
  or g45877 (n_16544, n_21982, wc163);
  not gc163 (wc163, n_16146);
  nand g45878 (n_16631, n_21942, n_23263);
  or g45879 (n_21900, n_16122, n_16420);
  nand g45880 (n_16605, n_21981, n_23266);
  or g45881 (n_21906, n_16125, n_16420);
  nand g45883 (n_24377, n_16671, n_16687);
  or g45884 (n_24378, n_16671, n_16687);
  nand g45885 (n_16688, n_24377, n_24378);
  or g45886 (n_21950, \data_stack_mem[7] [6], wc164);
  not gc164 (wc164, n_16633);
  or g45887 (n_21951, wc165, n_16633);
  not gc165 (wc165, \data_stack_mem[7] [6]);
  or g45888 (n_21876, n_16110, n_16420);
  or g45889 (n_22009, \data_stack_mem[6] [7], wc166);
  not gc166 (wc166, n_16668);
  or g45890 (n_16696, n_17317, wc167);
  not gc167 (wc167, n_21976);
  nand g45891 (n_16566, n_22017, n_22018);
  nand g45892 (n_21982, n_17423, n_21981);
  or g45893 (n_16744, n_17326, wc168);
  not gc168 (wc168, n_21967);
  or g45896 (n_16509, n_21943, wc169);
  not gc169 (wc169, n_16146);
  nand g45897 (n_22043, n_17694, n_16472);
  or g45898 (n_22012, \data_stack_mem[6] [7], n_16721);
  nand g45899 (n_22029, \data_stack_mem[7] [6], n_16625);
  nand g45900 (n_23263, n_16530, n_17388);
  or g45901 (n_22023, \data_stack_mem[9] [5], wc170);
  not gc170 (wc170, n_16532);
  nand g45902 (n_24379, n_16608, n_16622);
  or g45903 (n_24380, n_16608, n_16622);
  nand g45904 (n_16623, n_24379, n_24380);
  nand g45905 (n_23266, n_16564, n_17423);
  nand g45906 (n_16633, n_21846, n_23251);
  or g45907 (n_21987, n_16601, n_16625);
  nand g45910 (n_16668, n_21930, n_23257);
  nand g45911 (n_22005, n_22002, n_22003);
  nand g45912 (n_24381, n_16704, n_16802);
  or g45913 (n_24382, n_16704, n_16802);
  nand g45914 (n_16803, n_24381, n_24382);
  or g45916 (n_21871, n_21869, n_21870);
  nand g45917 (n_22004, n_17697, n_16493);
  nand g45918 (n_24383, n_16817, n_16820);
  or g45919 (n_24384, n_16817, n_16820);
  nand g45920 (n_16821, n_24383, n_24384);
  nand g45921 (n_17317, n_16154, n_21856);
  nand g45922 (n_16705, n_16704, n_21964);
  nand g45923 (n_24385, n_16511, n_16529);
  or g45924 (n_24386, n_16511, n_16529);
  nand g45925 (n_16530, n_24385, n_24386);
  nand g45926 (n_23251, n_16529, n_17464);
  nand g45927 (n_16721, n_21924, n_23254);
  nand g45928 (n_23257, n_16648, n_17449);
  nand g45929 (n_16625, n_21936, n_23260);
  nand g45930 (n_16532, n_21972, n_21973);
  nand g45932 (n_21981, \data_stack_mem[8] [5], n_16543);
  nand g45933 (n_24387, n_16546, n_16563);
  or g45934 (n_24388, n_16546, n_16563);
  nand g45935 (n_16564, n_24387, n_24388);
  nand g45936 (n_21976, n_16687, n_17465);
  nand g45937 (n_17694, n_21957, n_21958);
  nand g45938 (n_21931, n_17449, n_21930);
  nand g45939 (n_22017, n_17441, n_16472);
  nand g45940 (n_17326, n_16154, n_21859);
  nand g45941 (n_17693, n_17441, n_21991);
  nand g45943 (n_21943, n_17388, n_21942);
  nand g45944 (n_16342, n_21696, n_21697);
  nand g45945 (n_16344, n_21702, n_21703);
  nand g45946 (n_22018, \data_stack_mem[9] [4], n_16470);
  nand g45947 (n_16346, n_21708, n_21709);
  or g45948 (n_21930, \data_stack_mem[6] [6], wc171);
  not gc171 (wc171, n_16634);
  or g45949 (n_21859, \data_stack_mem[5] [7], n_16723);
  nand g45950 (n_16350, n_21720, n_21721);
  nand g45951 (n_24389, n_16673, n_16686);
  or g45952 (n_24390, n_16673, n_16686);
  nand g45953 (n_16687, n_24389, n_24390);
  nand g45954 (n_16340, n_21690, n_21691);
  nand g45955 (n_16338, n_21684, n_21685);
  nand g45956 (n_21972, n_17321, n_16493);
  nand g45957 (n_16336, n_21678, n_21679);
  nand g45958 (n_23254, n_16622, n_17466);
  nand g45959 (n_21964, n_16703, n_16697);
  or g45960 (n_21856, \data_stack_mem[5] [7], wc172);
  not gc172 (wc172, n_16670);
  or g45961 (n_21870, wc173, n_16419);
  not gc173 (wc173, n_16416);
  nand g45962 (n_21925, n_17466, n_21924);
  nand g45963 (n_24391, n_17382, n_16528);
  or g45964 (n_24392, n_17382, n_16528);
  nand g45965 (n_16529, n_24391, n_24392);
  nand g45966 (n_24393, n_16726, n_16734);
  or g45967 (n_24394, n_16726, n_16734);
  nand g45968 (n_16735, n_24393, n_24394);
  or g45969 (n_16801, n_21862, wc174);
  not gc174 (wc174, n_16697);
  nand g45971 (n_24395, n_16745, n_16750);
  or g45972 (n_24396, n_16745, n_16750);
  nand g45973 (n_16751, n_24395, n_24396);
  nand g45974 (n_17697, n_21852, n_21853);
  nand g45976 (n_16543, n_21771, n_23239);
  nand g45977 (n_24397, n_16637, n_16647);
  or g45978 (n_24398, n_16637, n_16647);
  nand g45979 (n_16648, n_24397, n_24398);
  nand g45980 (n_17696, n_17321, n_21961);
  nand g45981 (n_23260, n_16563, n_17460);
  or g45982 (n_21957, wc175, n_16470);
  not gc175 (wc175, \data_stack_mem[9] [4]);
  or g45983 (n_21958, wc176, n_16471);
  not gc176 (wc176, n_16470);
  or g45984 (n_21991, n_16429, wc177);
  not gc177 (wc177, n_16470);
  or g45985 (n_22042, n_16145, n_16470);
  or g45986 (n_21942, \data_stack_mem[8] [5], wc178);
  not gc178 (wc178, n_16508);
  nand g45987 (n_16348, n_21714, n_21715);
  nand g45988 (n_16508, n_21726, n_23233);
  or g45989 (n_21714, n_16128, n_16335);
  or g45990 (n_21720, n_16131, n_16335);
  or g45991 (n_16745, n_17345, wc179);
  not gc179 (wc179, n_21817);
  nand g45992 (n_16723, n_21783, n_23245);
  or g45993 (n_22003, n_16145, n_16492);
  nand g45994 (n_16634, n_21732, n_23236);
  nand g45995 (n_21847, n_17464, n_21846);
  or g45996 (n_16637, n_21790, wc180);
  not gc180 (wc180, n_16154);
  or g45997 (n_21973, \data_stack_mem[9] [4], wc181);
  not gc181 (wc181, n_16492);
  nand g45998 (n_21937, n_17460, n_21936);
  nand g45999 (n_16670, n_21789, n_23248);
  nand g46000 (n_21924, \data_stack_mem[6] [6], n_16607);
  or g46001 (n_21852, \data_stack_mem[9] [4], n_16492);
  nand g46003 (n_21869, n_17700, n_16393);
  or g46004 (n_16416, n_21805, n_16176);
  or g46005 (n_21678, n_16110, n_16335);
  or g46006 (n_21684, n_16113, n_16335);
  nand g46007 (n_24399, n_16548, n_16562);
  or g46008 (n_24400, n_16548, n_16562);
  nand g46009 (n_16563, n_24399, n_24400);
  or g46010 (n_21853, n_16429, wc182);
  not gc182 (wc182, n_16492);
  nand g46011 (n_23239, n_17315, n_16469);
  or g46012 (n_21690, n_16335, n_16116);
  or g46014 (n_21696, n_16119, n_16335);
  nand g46015 (n_24401, n_16449, n_16469);
  or g46016 (n_24402, n_16449, n_16469);
  nand g46017 (n_16470, n_24401, n_24402);
  nand g46018 (n_24403, n_16610, n_16621);
  or g46019 (n_24404, n_16610, n_16621);
  nand g46020 (n_16622, n_24403, n_24404);
  or g46022 (n_21702, n_16122, n_16335);
  or g46023 (n_21708, n_16125, n_16335);
  nand g46024 (n_23233, n_17316, n_16491);
  nand g46027 (n_24405, n_16475, n_16491);
  or g46028 (n_24406, n_16475, n_16491);
  nand g46029 (n_16492, n_24405, n_24406);
  or g46030 (n_21846, \data_stack_mem[7] [5], wc183);
  not gc183 (wc183, n_16510);
  nand g46031 (n_21790, n_17320, n_21789);
  nand g46032 (n_23248, n_16647, n_17320);
  nand g46033 (n_16607, n_21777, n_23242);
  nand g46034 (n_21733, n_17501, n_21732);
  nand g46035 (n_24407, n_16800, n_16702);
  or g46036 (n_24408, n_16800, n_16702);
  nand g46037 (n_16802, n_24407, n_24408);
  nand g46040 (n_16820, n_16819, n_16818);
  nand g46041 (n_21936, \data_stack_mem[7] [5], n_16545);
  or g46042 (n_16393, n_21748, n_16175);
  nand g46043 (n_17345, n_16156, n_21760);
  or g46044 (n_16610, n_21784, wc184);
  not gc184 (wc184, n_16154);
  nand g46045 (n_21841, n_16686, n_17329);
  nand g46046 (n_23245, n_16621, n_17330);
  nand g46047 (n_23236, n_16528, n_17501);
  nand g46050 (n_16703, n_16702, n_21808);
  nand g46052 (n_17335, n_16156, n_21757);
  nand g46053 (n_24411, n_16612, n_16620);
  or g46054 (n_24412, n_16612, n_16620);
  nand g46055 (n_16621, n_24411, n_24412);
  nand g46056 (n_16491, n_21765, n_21766);
  nand g46057 (n_21778, n_17332, n_21777);
  nand g46058 (n_16545, n_21837, n_21838);
  nand g46060 (n_21808, n_16700, n_16701);
  or g46061 (n_21789, \data_stack_mem[5] [6], wc185);
  not gc185 (wc185, n_16636);
  nand g46062 (n_23242, n_16562, n_17332);
  nand g46063 (n_21784, n_17330, n_21783);
  nand g46064 (n_24413, n_16514, n_16527);
  or g46065 (n_24414, n_16514, n_16527);
  nand g46066 (n_16528, n_24413, n_24414);
  nand g46067 (n_24415, n_16728, n_16733);
  or g46068 (n_24416, n_16728, n_16733);
  nand g46069 (n_16734, n_24415, n_24416);
  or g46070 (n_21732, \data_stack_mem[6] [5], wc186);
  not gc186 (wc186, n_16512);
  nand g46071 (n_24417, n_16746, n_16749);
  or g46072 (n_24418, n_16746, n_16749);
  nand g46073 (n_16750, n_24417, n_24418);
  or g46074 (n_21760, \data_stack_mem[4] [7], n_16725);
  nand g46075 (n_24419, n_16675, n_16685);
  or g46076 (n_24420, n_16675, n_16685);
  nand g46077 (n_16686, n_24419, n_24420);
  nand g46079 (n_16510, n_21648, n_23230);
  nand g46080 (n_24421, n_16639, n_16646);
  or g46081 (n_24422, n_16639, n_16646);
  nand g46082 (n_16647, n_24421, n_24422);
  nand g46083 (n_21804, n_21801, n_21802);
  nand g46084 (n_21832, n_21829, n_21830);
  nand g46085 (n_16472, n_21813, n_21814);
  or g46086 (n_21673, n_21671, n_21672);
  or g46087 (n_16475, n_21727, wc187);
  not gc187 (wc187, n_16146);
  or g46088 (n_21757, \data_stack_mem[4] [7], wc188);
  not gc188 (wc188, n_16672);
  or g46089 (n_21829, n_16444, n_17445);
  or g46090 (n_21830, n_21828, wc189);
  not gc189 (wc189, n_16468);
  nand g46091 (n_21777, \data_stack_mem[6] [5], n_16547);
  nand g46092 (n_21727, n_17316, n_21726);
  nand g46093 (n_21837, \data_stack_mem[7] [4], n_17445);
  or g46094 (n_16701, n_17359, wc190);
  not gc190 (wc190, n_21664);
  or g46095 (n_21672, wc191, n_16334);
  not gc191 (wc191, n_16331);
  nand g46096 (n_16493, n_21753, n_21754);
  or g46097 (n_16612, n_21637, wc192);
  not gc192 (wc192, n_16156);
  nand g46098 (n_16725, n_21636, n_23224);
  nand g46099 (n_21813, n_17325, n_16415);
  nand g46100 (n_21783, \data_stack_mem[5] [6], n_16609);
  or g46101 (n_16449, n_21772, wc193);
  not gc193 (wc193, n_16146);
  nand g46102 (n_21803, n_17699, n_16414);
  or g46104 (n_21802, n_17325, n_16415);
  nand g46105 (n_16636, n_21630, n_23221);
  or g46106 (n_21765, n_16489, wc194);
  not gc194 (wc194, n_17671);
  nand g46107 (n_16672, n_21642, n_23227);
  nand g46108 (n_24423, n_16550, n_16561);
  or g46109 (n_24424, n_16550, n_16561);
  nand g46110 (n_16562, n_24423, n_24424);
  or g46111 (n_16514, n_21631, wc195);
  not gc195 (wc195, n_16154);
  or g46112 (n_21766, wc196, n_17671);
  not gc196 (wc196, n_16489);
  nand g46114 (n_21747, n_21744, n_21745);
  or g46115 (n_16639, n_21643, wc197);
  not gc197 (wc197, n_16156);
  nand g46116 (n_16512, n_21555, n_23215);
  nand g46117 (n_23230, n_16489, n_17323);
  nand g46118 (n_21831, n_17644, n_16466);
  or g46119 (n_21661, wc198, n_16733);
  not gc198 (wc198, n_17362);
  nand g46120 (n_21643, n_17337, n_21642);
  or g46121 (n_21745, n_17324, n_16392);
  nand g46122 (n_21631, n_17331, n_21630);
  nand g46123 (n_23227, n_16646, n_17337);
  nand g46124 (n_24425, n_16477, n_16488);
  or g46125 (n_24426, n_16477, n_16488);
  nand g46126 (n_16489, n_24425, n_24426);
  nand g46127 (n_17448, n_16158, n_21601);
  nand g46128 (n_16609, n_21624, n_23218);
  nand g46129 (n_17359, n_16158, n_21598);
  nand g46130 (n_17698, n_16145, n_21652);
  nand g46131 (n_23221, n_16527, n_17331);
  nand g46132 (n_21772, n_17315, n_21771);
  nand g46133 (n_21814, \data_stack_mem[9] [3], n_16414);
  nand g46134 (n_21637, n_17413, n_21636);
  nand g46135 (n_17699, n_21657, n_21658);
  nand g46136 (n_21753, n_17324, n_16392);
  nand g46137 (n_23224, n_16620, n_17413);
  or g46138 (n_16331, n_21595, n_16176);
  nand g46139 (n_21664, n_16685, n_17349);
  or g46140 (n_16550, n_21625, wc199);
  not gc199 (wc199, n_16154);
  or g46141 (n_21726, \data_stack_mem[8] [4], wc200);
  not gc200 (wc200, n_16474);
  nand g46142 (n_21838, n_16466, n_16468);
  or g46143 (n_21828, n_16466, n_16467);
  nand g46144 (n_16547, n_21549, n_23212);
  nand g46145 (n_23215, n_17340, n_16488);
  nand g46146 (n_21671, n_17705, n_16308);
  nand g46147 (n_24427, n_16614, n_16619);
  or g46148 (n_24428, n_16614, n_16619);
  nand g46149 (n_16620, n_24427, n_24428);
  or g46152 (n_21642, \data_stack_mem[4] [6], wc201);
  not gc201 (wc201, n_16638);
  nand g46153 (n_21746, n_17702, n_16390);
  nand g46154 (n_16474, n_21471, n_23191);
  nand g46155 (n_24429, n_17410, n_16487);
  or g46156 (n_24430, n_17410, n_16487);
  nand g46157 (n_16488, n_24429, n_24430);
  nand g46158 (n_24431, n_16451, n_16465);
  or g46159 (n_24432, n_16451, n_16465);
  nand g46160 (n_16466, n_24431, n_24432);
  or g46162 (n_21657, n_16351, n_16415);
  nand g46163 (n_21625, n_17339, n_21624);
  nand g46164 (n_17671, n_21570, n_21571);
  nand g46165 (n_21771, \data_stack_mem[8] [4], n_16448);
  nand g46166 (n_24433, n_16395, n_16413);
  or g46167 (n_24434, n_16395, n_16413);
  nand g46168 (n_16414, n_24433, n_24434);
  or g46169 (n_21754, \data_stack_mem[9] [3], wc202);
  not gc202 (wc202, n_16390);
  nand g46170 (n_21652, \data_stack_mem[9] [3], n_16415);
  or g46171 (n_21630, \data_stack_mem[5] [5], wc203);
  not gc203 (wc203, n_16513);
  nand g46172 (n_23212, n_16465, n_17338);
  nand g46173 (n_24435, n_16516, n_16526);
  or g46174 (n_24436, n_16516, n_16526);
  nand g46175 (n_16527, n_24435, n_24436);
  or g46176 (n_21744, n_16390, wc204);
  not gc204 (wc204, n_17701);
  nand g46177 (n_24437, n_16641, n_16645);
  or g46178 (n_24438, n_16641, n_16645);
  nand g46179 (n_16646, n_24437, n_24438);
  or g46180 (n_21601, \data_stack_mem[3] [7], n_16727);
  nand g46181 (n_21636, \data_stack_mem[4] [6], n_16611);
  or g46182 (n_21598, \data_stack_mem[3] [7], wc205);
  not gc205 (wc205, n_16674);
  nand g46183 (n_23218, n_16561, n_17339);
  or g46185 (n_21571, n_16444, wc206);
  not gc206 (wc206, n_16490);
  nand g46186 (n_16513, n_21429, n_23182);
  nand g46187 (n_24439, n_16747, n_16748);
  or g46188 (n_24440, n_16747, n_16748);
  nand g46189 (n_16749, n_24439, n_24440);
  nand g46191 (n_24441, n_16371, n_16389);
  or g46192 (n_24442, n_16371, n_16389);
  nand g46193 (n_16390, n_24441, n_24442);
  nand g46194 (n_16349, n_21423, n_21424);
  nand g46195 (n_21565, n_21563, n_21564);
  nand g46196 (n_16674, n_21489, n_23200);
  or g46197 (n_16395, n_21544, wc207);
  not gc207 (wc207, n_16146);
  nand g46198 (n_17701, n_16145, n_21574);
  nand g46199 (n_24443, n_16453, n_16464);
  or g46200 (n_24444, n_16453, n_16464);
  nand g46201 (n_16465, n_24443, n_24444);
  nand g46202 (n_23191, n_17333, n_16389);
  nand g46203 (n_21624, \data_stack_mem[5] [5], n_16549);
  nand g46204 (n_16347, n_21417, n_21418);
  nand g46205 (n_21556, n_17340, n_21555);
  nand g46206 (n_21594, n_21591, n_21592);
  nand g46207 (n_17702, n_21579, n_21580);
  nand g46208 (n_16345, n_21411, n_21412);
  or g46209 (n_16308, n_21517, n_16175);
  nand g46212 (n_16343, n_21405, n_21406);
  nand g46213 (n_16337, n_21387, n_21388);
  nand g46214 (n_16341, n_21399, n_21400);
  or g46215 (n_16516, n_21496, wc208);
  not gc208 (wc208, n_16156);
  nand g46216 (n_24445, n_16552, n_16560);
  or g46217 (n_24446, n_16552, n_16560);
  nand g46218 (n_16561, n_24445, n_24446);
  nand g46219 (n_16727, n_21483, n_23197);
  nand g46220 (n_16611, n_21477, n_23194);
  nand g46221 (n_16339, n_21393, n_21394);
  or g46222 (n_21648, \data_stack_mem[7] [4], wc209);
  not gc209 (wc209, n_16490);
  or g46223 (n_17410, n_21430, wc210);
  not gc210 (wc210, n_16154);
  nand g46224 (n_16733, n_21612, n_21613);
  nand g46225 (n_16638, n_21495, n_23203);
  nand g46226 (n_16415, n_21618, n_21619);
  nand g46227 (n_16448, n_21543, n_23209);
  nand g46228 (n_16263, n_21381, n_21382);
  or g46229 (n_21570, n_16467, n_16490);
  or g46230 (n_16747, n_16730, wc211);
  not gc211 (wc211, n_21520);
  or g46231 (n_16552, n_21478, wc212);
  not gc212 (wc212, n_16156);
  or g46232 (n_21563, \data_stack_mem[7] [4], n_16468);
  nand g46233 (n_16389, n_21525, n_21526);
  nand g46234 (n_21564, \data_stack_mem[7] [4], n_16468);
  nand g46235 (n_21544, n_17334, n_21543);
  or g46236 (n_24447, wc213, n_16699);
  not gc213 (wc213, n_16698);
  or g46237 (n_24448, n_16698, wc214);
  not gc214 (wc214, n_16699);
  nand g46238 (n_16700, n_24447, n_24448);
  or g46239 (n_21555, \data_stack_mem[6] [4], wc215);
  not gc215 (wc215, n_16476);
  or g46240 (n_21592, n_17343, n_16330);
  nand g46241 (n_21550, n_17338, n_21549);
  nand g46242 (n_21484, n_17377, n_21483);
  nand g46244 (n_16549, n_21465, n_23188);
  nand g46245 (n_16685, n_21531, n_21532);
  nand g46246 (n_23197, n_17377, n_16619);
  nand g46247 (n_23194, n_16560, n_17364);
  nand g46248 (n_21430, n_17508, n_21429);
  nand g46249 (n_21496, n_17352, n_21495);
  nand g46250 (n_23203, n_16526, n_17352);
  or g46251 (n_21612, wc216, n_16732);
  not gc216 (wc216, n_17687);
  nand g46252 (n_21618, n_17343, n_16330);
  or g46253 (n_21613, n_17687, wc217);
  not gc217 (wc217, n_16732);
  nand g46254 (n_23200, n_17418, n_16645);
  nand g46255 (n_21490, n_17418, n_21489);
  or g46256 (n_21423, n_16131, n_16262);
  nand g46257 (n_23182, n_16487, n_17508);
  or g46258 (n_21417, n_16128, n_16262);
  or g46259 (n_21411, n_16125, n_16262);
  or g46260 (n_21405, n_16122, n_16262);
  or g46261 (n_21399, n_16119, n_16262);
  or g46262 (n_21393, n_16262, n_16116);
  or g46263 (n_16453, n_21466, wc218);
  not gc218 (wc218, n_16154);
  nand g46264 (n_16490, n_21441, n_23185);
  nand g46265 (n_16800, n_16699, n_16698);
  or g46266 (n_21579, n_16391, n_16392);
  or g46267 (n_21580, n_16351, wc219);
  not gc219 (wc219, n_16392);
  or g46268 (n_16371, n_21472, wc220);
  not gc220 (wc220, n_16146);
  or g46269 (n_21381, n_16110, n_16262);
  or g46270 (n_21387, n_16113, n_16262);
  or g46271 (n_21574, \data_stack_mem[9] [3], wc221);
  not gc221 (wc221, n_16392);
  nand g46272 (n_23209, n_17334, n_16413);
  nand g46273 (n_16730, n_16160, n_21451);
  or g46274 (n_21520, wc222, n_16732);
  not gc222 (wc222, n_17374);
  nand g46275 (n_24449, n_16554, n_16559);
  or g46276 (n_24450, n_16554, n_16559);
  nand g46277 (n_16560, n_24449, n_24450);
  nand g46278 (n_16413, n_21606, n_21607);
  nand g46279 (n_21472, n_17333, n_21471);
  nand g46280 (n_23185, n_16387, n_17341);
  nand g46281 (n_24451, n_17346, n_16486);
  or g46282 (n_24452, n_17346, n_16486);
  nand g46283 (n_16487, n_24451, n_24452);
  or g46284 (n_21489, \data_stack_mem[3] [6], wc223);
  not gc223 (wc223, n_16640);
  nand g46285 (n_17687, n_21447, n_21448);
  or g46286 (n_21495, \data_stack_mem[4] [5], wc224);
  not gc224 (wc224, n_16515);
  nand g46287 (n_21619, \data_stack_mem[9] [2], n_16329);
  nand g46288 (n_16392, n_21537, n_21538);
  or g46289 (n_21429, \data_stack_mem[5] [4], wc225);
  not gc225 (wc225, n_16478);
  nand g46290 (n_24453, n_16518, n_16525);
  or g46291 (n_24454, n_16518, n_16525);
  nand g46292 (n_16526, n_24453, n_24454);
  nand g46293 (n_23188, n_16464, n_17363);
  or g46294 (n_21531, wc226, n_16684);
  not gc226 (wc226, n_17691);
  or g46295 (n_21532, n_17691, wc227);
  not gc227 (wc227, n_16684);
  nand g46296 (n_21483, \data_stack_mem[3] [6], n_16613);
  nand g46297 (n_21516, n_21513, n_21514);
  nand g46298 (n_21593, n_17704, n_16329);
  nand g46299 (n_21549, \data_stack_mem[6] [4], n_16450);
  or g46300 (n_21591, n_16329, wc228);
  not gc228 (wc228, n_17703);
  nand g46301 (n_16476, n_21285, n_23164);
  nand g46303 (n_21543, \data_stack_mem[8] [3], n_16394);
  nand g46304 (n_16468, n_21501, n_23206);
  or g46305 (n_16698, n_16679, wc229);
  not gc229 (wc229, n_21454);
  nand g46306 (n_21478, n_17364, n_21477);
  or g46307 (n_21526, wc230, n_17676);
  not gc230 (wc230, n_16387);
  or g46308 (n_21525, n_16387, wc231);
  not gc231 (wc231, n_17676);
  nand g46309 (n_21466, n_17363, n_21465);
  or g46310 (n_17346, n_21310, wc232);
  not gc232 (wc232, n_16156);
  or g46311 (n_21447, n_16676, n_16729);
  or g46312 (n_21448, n_16677, wc233);
  not gc233 (wc233, n_16729);
  nand g46314 (n_16619, n_21459, n_21460);
  nand g46315 (n_21537, n_17344, n_16307);
  nand g46316 (n_16515, n_21309, n_23176);
  nand g46317 (n_21477, \data_stack_mem[4] [5], n_16551);
  nand g46318 (n_17691, n_21327, n_21328);
  nand g46319 (n_21465, \data_stack_mem[5] [4], n_16452);
  nand g46320 (n_16679, n_16160, n_21340);
  nand g46321 (n_24455, n_16373, n_16386);
  or g46322 (n_24456, n_16373, n_16386);
  nand g46323 (n_16387, n_24455, n_24456);
  nand g46324 (n_21454, n_17360, n_16684);
  or g46325 (n_21471, \data_stack_mem[8] [3], wc234);
  not gc234 (wc234, n_16370);
  nand g46326 (n_23206, n_16411, n_17342);
  nand g46328 (n_16450, n_21291, n_23167);
  nand g46329 (n_24457, n_16310, n_16328);
  or g46330 (n_24458, n_16310, n_16328);
  nand g46331 (n_16329, n_24457, n_24458);
  or g46332 (n_21514, n_17344, n_16307);
  nand g46333 (n_16613, n_21297, n_23170);
  or g46334 (n_21451, \data_stack_mem[2] [7], n_16729);
  nand g46335 (n_16640, n_21303, n_23173);
  or g46336 (n_21607, wc235, n_17664);
  not gc235 (wc235, n_16411);
  nand g46337 (n_24459, n_16455, n_16463);
  or g46338 (n_24460, n_16455, n_16463);
  nand g46339 (n_16464, n_24459, n_24460);
  or g46340 (n_21606, n_16411, wc236);
  not gc236 (wc236, n_17664);
  nand g46341 (n_23164, n_16386, n_17351);
  or g46342 (n_21376, n_21374, n_21375);
  nand g46343 (n_16394, n_21279, n_23161);
  nand g46344 (n_16478, n_21225, n_23149);
  nand g46345 (n_17676, n_21315, n_21316);
  or g46346 (n_21460, n_17684, wc237);
  not gc237 (wc237, n_16618);
  or g46347 (n_21459, wc238, n_16618);
  not gc238 (wc238, n_17684);
  nand g46348 (n_23161, n_17357, n_16328);
  or g46349 (n_21375, wc239, n_16261);
  not gc239 (wc239, n_16258);
  nand g46350 (n_17703, n_16145, n_21331);
  or g46351 (n_16455, n_21274, wc240);
  not gc240 (wc240, n_16156);
  nand g46352 (n_17704, n_21336, n_21337);
  or g46353 (n_21513, n_16305, wc241);
  not gc241 (wc241, n_17707);
  nand g46354 (n_16551, n_21273, n_23158);
  nand g46355 (n_21515, n_17708, n_16305);
  or g46356 (n_21340, \data_stack_mem[2] [7], wc242);
  not gc242 (wc242, n_16678);
  nand g46357 (n_24461, n_16375, n_16385);
  or g46358 (n_24462, n_16375, n_16385);
  nand g46359 (n_16386, n_24461, n_24462);
  nand g46360 (n_23167, n_16410, n_17355);
  or g46361 (n_16310, n_21280, wc243);
  not gc243 (wc243, n_16146);
  nand g46362 (n_21298, n_17402, n_21297);
  nand g46363 (n_23149, n_17379, n_16385);
  nand g46364 (n_23170, n_16559, n_17402);
  or g46366 (n_21538, \data_stack_mem[9] [2], wc244);
  not gc244 (wc244, n_16305);
  nand g46367 (n_21310, n_17510, n_21309);
  nand g46368 (n_23173, n_16525, n_17375);
  nand g46369 (n_16645, n_21360, n_21361);
  nand g46370 (n_24463, n_16397, n_16410);
  or g46371 (n_24464, n_16397, n_16410);
  nand g46372 (n_16411, n_24463, n_24464);
  nand g46373 (n_16452, n_21231, n_23152);
  nand g46374 (n_16370, n_21219, n_23146);
  nand g46375 (n_17664, n_21435, n_21436);
  or g46376 (n_21327, n_16677, n_16678);
  or g46377 (n_21328, n_16676, wc245);
  not gc245 (wc245, n_16678);
  nand g46378 (n_23176, n_16486, n_17510);
  nand g46379 (n_16729, n_21321, n_23179);
  nand g46380 (n_21304, n_17375, n_21303);
  or g46381 (n_21336, n_16264, n_16330);
  nand g46384 (n_21501, \data_stack_mem[7] [3], n_16412);
  or g46385 (n_21435, n_16353, n_16412);
  or g46386 (n_21303, \data_stack_mem[3] [5], wc246);
  not gc246 (wc246, n_16517);
  nand g46387 (n_24465, n_17419, n_16384);
  or g46388 (n_24466, n_17419, n_16384);
  nand g46389 (n_16385, n_24465, n_24466);
  nand g46390 (n_21297, \data_stack_mem[3] [5], n_16553);
  nand g46392 (n_21331, \data_stack_mem[9] [2], n_16330);
  nand g46393 (n_24467, n_16284, n_16304);
  or g46394 (n_24468, n_16284, n_16304);
  nand g46395 (n_16305, n_24467, n_24468);
  or g46396 (n_21316, n_16353, wc247);
  not gc247 (wc247, n_16388);
  or g46397 (n_16258, n_21262, n_16176);
  or g46398 (n_21361, n_17686, wc248);
  not gc248 (wc248, n_16644);
  nand g46399 (n_23179, n_17319, n_16618);
  nand g46400 (n_24469, n_16399, n_16409);
  or g46401 (n_24470, n_16399, n_16409);
  nand g46402 (n_16410, n_24469, n_24470);
  or g46403 (n_21360, wc249, n_16644);
  not gc249 (wc249, n_17686);
  nand g46404 (n_23146, n_17358, n_16304);
  or g46405 (n_21315, n_17260, n_16388);
  nand g46406 (n_17684, n_21237, n_21238);
  nand g46407 (n_21280, n_17357, n_21279);
  nand g46408 (n_16678, n_21243, n_23155);
  or g46409 (n_21441, \data_stack_mem[7] [3], wc250);
  not gc250 (wc250, n_16388);
  nand g46410 (n_23158, n_16463, n_17452);
  or g46412 (n_21309, \data_stack_mem[4] [4], wc251);
  not gc251 (wc251, n_16479);
  nand g46413 (n_23152, n_16409, n_17380);
  nand g46414 (n_21274, n_17452, n_21273);
  nand g46415 (n_21286, n_17351, n_21285);
  or g46416 (n_16375, n_21226, wc252);
  not gc252 (wc252, n_16154);
  nand g46417 (n_24471, n_16481, n_16485);
  or g46418 (n_24472, n_16481, n_16485);
  nand g46419 (n_16486, n_24471, n_24472);
  nand g46420 (n_24473, n_16457, n_16462);
  or g46421 (n_24474, n_16457, n_16462);
  nand g46422 (n_16463, n_24473, n_24474);
  nand g46423 (n_17707, n_16145, n_21247);
  or g46424 (n_17419, n_21049, wc253);
  not gc253 (wc253, n_16156);
  nand g46425 (n_21279, \data_stack_mem[8] [2], n_16309);
  nand g46426 (n_21355, n_21352, n_21353);
  nand g46427 (n_16517, n_21177, n_23137);
  or g46428 (n_21285, \data_stack_mem[6] [3], wc254);
  not gc254 (wc254, n_16372);
  nand g46429 (n_24475, n_16401, n_16408);
  or g46430 (n_24476, n_16401, n_16408);
  nand g46431 (n_16409, n_24475, n_24476);
  nand g46432 (n_16304, n_21267, n_21268);
  nand g46433 (n_17686, n_21204, n_21205);
  nand g46434 (n_21273, \data_stack_mem[4] [4], n_16454);
  nand g46435 (n_21321, \data_stack_mem[2] [6], n_16615);
  nand g46436 (n_24477, n_16556, n_16558);
  or g46437 (n_24478, n_16556, n_16558);
  nand g46438 (n_16559, n_24477, n_24478);
  nand g46439 (n_16330, n_21060, n_23125);
  nand g46440 (n_16388, n_21198, n_23143);
  nand g46441 (n_16479, n_21048, n_23122);
  nand g46442 (n_16412, n_21366, n_21367);
  or g46443 (n_21238, n_16616, wc255);
  not gc255 (wc255, n_16615);
  nand g46444 (n_21374, n_17711, n_16237);
  nand g46445 (n_23155, n_17322, n_16644);
  nand g46447 (n_21292, n_17355, n_21291);
  nand g46448 (n_21226, n_17379, n_21225);
  nand g46449 (n_16553, n_21171, n_23134);
  or g46450 (n_21237, n_16593, n_16615);
  or g46451 (n_16284, n_21220, wc256);
  not gc256 (wc256, n_16146);
  or g46452 (n_16399, n_21232, wc257);
  not gc257 (wc257, n_16154);
  nand g46453 (n_21262, n_21260, n_21261);
  nand g46454 (n_17708, n_21252, n_21253);
  or g46456 (n_16237, n_21214, n_16175);
  or g46457 (n_21260, n_16257, n_17710);
  nand g46458 (n_21261, n_17710, n_16257);
  or g46459 (n_21225, \data_stack_mem[5] [3], wc258);
  not gc258 (wc258, n_16374);
  nand g46460 (n_23137, n_17457, n_16485);
  nand g46461 (n_21291, \data_stack_mem[6] [3], n_16396);
  nand g46462 (n_21232, n_17380, n_21231);
  nand g46463 (n_23143, n_16301, n_17446);
  or g46464 (n_16401, n_21166, wc259);
  not gc259 (wc259, n_16156);
  nand g46465 (n_16615, n_21183, n_23140);
  or g46466 (n_21247, \data_stack_mem[9] [2], wc260);
  not gc260 (wc260, n_16307);
  or g46467 (n_21253, n_16264, wc261);
  not gc261 (wc261, n_16307);
  or g46468 (n_21252, n_16306, n_16307);
  nand g46469 (n_24479, n_16520, n_16524);
  or g46470 (n_24480, n_16520, n_16524);
  nand g46471 (n_16525, n_24479, n_24480);
  or g46472 (n_21267, n_16301, wc262);
  not gc262 (wc262, n_17680);
  or g46473 (n_21268, wc263, n_17680);
  not gc263 (wc263, n_16301);
  nand g46475 (n_23122, n_16384, n_17507);
  nand g46476 (n_16309, n_20943, n_23095);
  nand g46477 (n_21049, n_17507, n_21048);
  nand g46478 (n_21178, n_17457, n_21177);
  nand g46479 (n_21354, n_17665, n_16326);
  nand g46480 (n_23125, n_16257, n_17370);
  or g46481 (n_21352, n_16279, n_17431);
  or g46482 (n_21204, n_16616, n_16642);
  or g46483 (n_21205, n_16593, wc264);
  not gc264 (wc264, n_16642);
  nand g46484 (n_16372, n_21030, n_23113);
  or g46485 (n_21243, \data_stack_mem[2] [6], wc265);
  not gc265 (wc265, n_16642);
  nand g46486 (n_21220, n_17358, n_21219);
  nand g46487 (n_21366, \data_stack_mem[7] [2], n_17431);
  nand g46488 (n_16454, n_21165, n_23131);
  or g46489 (n_21353, n_21351, wc266);
  not gc266 (wc266, n_16327);
  nand g46490 (n_23134, n_17395, n_16462);
  nand g46491 (n_24481, n_16239, n_16256);
  or g46492 (n_24482, n_16239, n_16256);
  nand g46493 (n_16257, n_24481, n_24482);
  nand g46494 (n_16188, n_21123, n_21124);
  nand g46495 (n_16190, n_21135, n_21136);
  nand g46496 (n_16462, n_21084, n_21085);
  nand g46497 (n_16189, n_21129, n_21130);
  nand g46498 (n_21184, n_17403, n_21183);
  nand g46499 (n_21367, n_16326, n_16327);
  or g46500 (n_21048, \data_stack_mem[4] [3], wc267);
  not gc267 (wc267, n_16376);
  nand g46501 (n_16192, n_21147, n_21148);
  or g46502 (n_21177, \data_stack_mem[3] [4], wc268);
  not gc268 (wc268, n_16480);
  nand g46503 (n_24483, n_16286, n_16300);
  or g46504 (n_24484, n_16286, n_16300);
  nand g46505 (n_16301, n_24483, n_24484);
  nand g46506 (n_23113, n_16300, n_17381);
  nand g46507 (n_23131, n_17400, n_16408);
  nand g46508 (n_21214, n_21212, n_21213);
  nand g46509 (n_16384, n_21078, n_21079);
  nand g46510 (n_21231, \data_stack_mem[5] [3], n_16398);
  nand g46511 (n_16187, n_21117, n_21118);
  or g46512 (n_21219, \data_stack_mem[8] [2], wc269);
  not gc269 (wc269, n_16283);
  nand g46513 (n_16194, n_21159, n_21160);
  nand g46515 (n_16642, n_21042, n_23119);
  nand g46516 (n_21166, n_17400, n_21165);
  or g46517 (n_16485, wc270, n_21019);
  not gc270 (wc270, n_21018);
  nand g46518 (n_16191, n_21141, n_21142);
  nand g46519 (n_21172, n_17395, n_21171);
  nand g46520 (n_23140, n_16558, n_17403);
  or g46521 (n_21351, n_16302, n_16326);
  nand g46523 (n_16193, n_21153, n_21154);
  nand g46524 (n_16307, n_21066, n_23128);
  nand g46525 (n_23095, n_17422, n_16256);
  nand g46526 (n_16396, n_21036, n_23116);
  nand g46527 (n_16374, n_20949, n_23098);
  nand g46528 (n_21043, n_17398, n_21042);
  nand g46529 (n_23116, n_16325, n_17376);
  nand g46530 (n_23128, n_16234, n_17372);
  or g46531 (n_21141, n_16122, n_16186);
  nand g46532 (n_23098, n_16299, n_17383);
  or g46533 (n_21135, n_16119, n_16186);
  or g46536 (n_21123, n_16113, n_16186);
  nand g46537 (n_21183, \data_stack_mem[2] [5], n_16555);
  or g46538 (n_21129, n_16186, n_16116);
  or g46541 (n_21159, n_16131, n_16186);
  nand g46542 (n_16408, n_21072, n_21073);
  nand g46543 (n_21085, n_16460, n_17672);
  nand g46544 (n_16283, n_20937, n_23092);
  nand g46545 (n_17680, n_21054, n_21055);
  or g46546 (n_21084, n_17672, n_16460);
  nand g46547 (n_21018, n_17669, n_16484);
  or g46548 (n_21212, n_16234, n_17713);
  nand g46549 (n_21165, \data_stack_mem[4] [3], n_16400);
  nand g46550 (n_23119, n_16524, n_17398);
  nand g46551 (n_16376, n_20868, n_23083);
  or g46552 (n_21117, n_16110, n_16186);
  or g46553 (n_21153, n_16128, n_16186);
  nand g46554 (n_24485, n_16312, n_16325);
  or g46555 (n_24486, n_16312, n_16325);
  nand g46556 (n_16326, n_24485, n_24486);
  nand g46557 (n_21213, n_17713, n_16234);
  nand g46558 (n_16480, n_20967, n_23107);
  or g46559 (n_21147, n_16125, n_16186);
  nand g46560 (n_21171, \data_stack_mem[3] [4], n_16456);
  nand g46561 (n_16398, n_20955, n_23101);
  nand g46562 (n_21193, n_21191, n_21192);
  nand g46563 (n_24487, n_16288, n_16299);
  or g46564 (n_24488, n_16288, n_16299);
  nand g46565 (n_16300, n_24487, n_24488);
  nand g46566 (n_21103, n_21100, n_21101);
  nand g46567 (n_24489, n_16290, n_16298);
  or g46568 (n_24490, n_16290, n_16298);
  nand g46569 (n_16299, n_24489, n_24490);
  or g46570 (n_21198, \data_stack_mem[7] [2], wc271);
  not gc271 (wc271, n_16303);
  nand g46571 (n_23092, n_17421, n_16233);
  or g46572 (n_16288, n_20950, wc272);
  not gc272 (wc272, n_16154);
  nand g46574 (n_23083, n_17327, n_16298);
  or g46575 (n_21042, \data_stack_mem[2] [5], wc273);
  not gc273 (wc273, n_16519);
  nand g46578 (n_21019, n_21016, n_21017);
  nand g46580 (n_16400, n_20874, n_23086);
  or g46582 (n_21054, n_16302, n_16303);
  nand g46583 (n_24491, n_16314, n_16324);
  or g46584 (n_24492, n_16314, n_16324);
  nand g46585 (n_16325, n_24491, n_24492);
  nand g46586 (n_23107, n_16381, n_17399);
  or g46587 (n_21055, n_16279, wc274);
  not gc274 (wc274, n_16303);
  or g46588 (n_21191, \data_stack_mem[7] [2], n_16327);
  nand g46589 (n_24493, n_16215, n_16233);
  or g46590 (n_24494, n_16215, n_16233);
  nand g46591 (n_16234, n_24493, n_24494);
  or g46592 (n_16186, n_16144, wc275);
  not gc275 (wc275, n_21112);
  nand g46593 (n_17657, n_20886, n_20887);
  nand g46594 (n_16555, n_20973, n_23110);
  nand g46595 (n_23101, n_16324, n_17386);
  nand g46596 (n_21192, \data_stack_mem[7] [2], n_16327);
  nand g46597 (n_21031, n_17381, n_21030);
  nand g46598 (n_16456, n_20961, n_23104);
  nand g46599 (n_20974, n_17350, n_20973);
  or g46600 (n_16290, n_20869, wc276);
  not gc276 (wc276, n_16156);
  or g46601 (n_21101, \data_stack_mem[7] [1], n_21099);
  nand g46602 (n_20950, n_17383, n_20949);
  or g46603 (n_16314, n_20956, wc277);
  not gc277 (wc277, n_16154);
  nand g46605 (n_17650, n_20880, n_20881);
  nand g46606 (n_20896, n_20894, n_20895);
  or g46607 (n_20967, \data_stack_mem[3] [3], wc278);
  not gc278 (wc278, n_16383);
  or g46608 (n_20886, n_16382, n_16383);
  or g46609 (n_20887, n_16364, wc279);
  not gc279 (wc279, n_16383);
  nand g46610 (n_16519, n_20931, n_20932);
  nand g46611 (n_23104, n_16406, n_17406);
  nand g46612 (n_16303, n_20910, n_23089);
  nand g46613 (n_16298, n_20862, n_20863);
  nand g46614 (n_24495, n_16316, n_16323);
  or g46615 (n_24496, n_16316, n_16323);
  nand g46616 (n_16324, n_24495, n_24496);
  nand g46617 (n_23086, n_17407, n_16323);
  nand g46618 (n_16233, n_21024, n_21025);
  nand g46620 (n_23110, n_17350, n_16460);
  or g46621 (n_21030, \data_stack_mem[6] [2], wc280);
  not gc280 (wc280, n_16285);
  nand g46622 (n_21037, n_17376, n_21036);
  nand g46623 (n_16327, n_21108, n_21109);
  or g46625 (n_21100, n_16210, n_17393);
  nand g46626 (n_16285, n_20796, n_23068);
  or g46627 (n_21099, n_21098, wc281);
  not gc281 (wc281, n_16169);
  nand g46628 (n_16383, n_20763, n_23065);
  nand g46629 (n_20956, n_17386, n_20955);
  or g46630 (n_21015, n_17404, wc282);
  not gc282 (wc282, n_16482);
  or g46632 (n_21016, n_21014, n_16482);
  nand g46633 (n_20869, n_17327, n_20868);
  nand g46634 (n_24497, n_16378, n_16380);
  or g46635 (n_24498, n_16378, n_16380);
  nand g46636 (n_16381, n_24497, n_24498);
  or g46637 (n_20895, \data_stack_mem[2] [4], wc283);
  not gc283 (wc283, n_16482);
  or g46638 (n_21025, wc284, n_17682);
  not gc284 (wc284, n_16231);
  or g46639 (n_21024, n_16231, wc285);
  not gc285 (wc285, n_17682);
  nand g46640 (n_21036, \data_stack_mem[6] [2], n_16311);
  or g46641 (n_20894, wc286, n_16482);
  not gc286 (wc286, \data_stack_mem[2] [4]);
  nand g46642 (n_20931, n_17404, n_16482);
  nand g46643 (n_23089, n_16231, n_17394);
  nand g46646 (n_16323, n_20925, n_20926);
  nand g46647 (n_20973, \data_stack_mem[2] [4], n_16461);
  or g46648 (n_20880, n_16364, n_16407);
  or g46649 (n_20881, n_16382, wc287);
  not gc287 (wc287, n_16407);
  or g46650 (n_16316, n_20875, wc288);
  not gc288 (wc288, n_16156);
  or g46652 (n_20949, \data_stack_mem[5] [2], wc289);
  not gc289 (wc289, n_16287);
  nand g46653 (n_20961, \data_stack_mem[3] [3], n_16407);
  nand g46654 (n_21108, \data_stack_mem[7] [1], n_17393);
  nand g46655 (n_24499, n_16403, n_16405);
  or g46656 (n_24500, n_16403, n_16405);
  nand g46657 (n_16406, n_24499, n_24500);
  nand g46658 (n_20875, n_17407, n_20874);
  nand g46659 (n_23068, n_16230, n_17397);
  nand g46660 (n_21102, n_17674, n_16255);
  or g46661 (n_21098, n_16255, n_16149);
  nand g46662 (n_23065, n_16295, n_17408);
  nand g46663 (n_16482, n_20808, n_23074);
  nand g46664 (n_17710, n_20979, n_20980);
  nand g46665 (n_19450, n_19448, n_19449);
  or g46666 (n_16215, n_20938, wc290);
  not gc290 (wc290, n_16146);
  or g46667 (n_20868, \data_stack_mem[4] [2], wc291);
  not gc291 (wc291, n_16289);
  or g46668 (n_16239, n_20944, wc292);
  not gc292 (wc292, n_16146);
  nand g46669 (n_16311, n_20802, n_23071);
  nand g46671 (n_24501, n_16217, n_16230);
  or g46672 (n_24502, n_16217, n_16230);
  nand g46673 (n_16231, n_24501, n_24502);
  nand g46674 (n_16699, n_17717, n_16162);
  nand g46675 (n_17713, n_20985, n_20986);
  nand g46677 (n_21001, n_20998, n_20999);
  nand g46678 (n_19438, n_19436, n_19437);
  nand g46680 (n_16407, n_20820, n_23080);
  nand g46681 (n_16461, n_20814, n_23077);
  nand g46682 (n_20955, \data_stack_mem[5] [2], n_16313);
  nand g46683 (n_16287, n_20745, n_23059);
  or g46685 (n_21109, n_16240, wc293);
  not gc293 (wc293, n_16255);
  nand g46686 (n_17653, n_20739, n_20740);
  or g46687 (n_20986, n_16195, wc294);
  not gc294 (wc294, n_16236);
  or g46688 (n_20985, n_16235, n_16236);
  nand g46689 (n_23074, n_17347, n_16380);
  nand g46690 (n_23080, n_16321, n_17414);
  or g46691 (n_20979, n_16172, n_16235);
  or g46692 (n_20980, wc295, n_16195);
  not gc295 (wc295, n_16172);
  nand g46693 (n_20874, \data_stack_mem[4] [2], n_16315);
  nand g46694 (n_20938, n_17421, n_20937);
  nand g46695 (n_20944, n_17422, n_20943);
  nand g46696 (n_24503, n_16242, n_16254);
  or g46697 (n_24504, n_16242, n_16254);
  nand g46698 (n_16255, n_24503, n_24504);
  nand g46699 (n_16313, n_20751, n_23062);
  nand g46700 (n_16748, n_23013, n_23014);
  nand g46702 (n_17642, n_20757, n_20758);
  or g46703 (n_20999, n_16172, wc296);
  not gc296 (wc296, n_16145);
  or g46705 (n_21060, wc297, n_16172);
  not gc297 (wc297, \data_stack_mem[9] [1]);
  nand g46706 (n_17717, n_17911, n_22999);
  nand g46707 (n_23077, n_17444, n_16405);
  nand g46708 (n_20815, n_17444, n_20814);
  nand g46709 (n_23059, n_16229, n_17405);
  nand g46710 (n_24505, n_16219, n_16229);
  or g46711 (n_24506, n_16219, n_16229);
  nand g46712 (n_16230, n_24505, n_24506);
  or g46714 (n_20739, n_16296, n_16297);
  or g46715 (n_20763, \data_stack_mem[3] [2], wc298);
  not gc298 (wc298, n_16297);
  or g46717 (n_21066, \data_stack_mem[9] [1], wc299);
  not gc299 (wc299, n_16236);
  nand g46718 (n_16289, n_20706, n_23047);
  nand g46719 (n_23071, n_16254, n_17328);
  or g46720 (n_20740, n_16268, wc300);
  not gc300 (wc300, n_16297);
  or g46721 (n_17689, n_20920, n_16178);
  nand g46722 (n_20809, n_17347, n_20808);
  or g46724 (n_17711, n_20857, n_16178);
  nand g46725 (n_16789, n_17750, n_16788);
  or g46726 (n_20943, wc301, n_16238);
  not gc301 (wc301, \data_stack_mem[8] [1]);
  nand g46727 (n_16185, n_17757, n_16184);
  nand g46728 (n_17682, n_20838, n_20839);
  nand g46729 (n_20830, n_20828, n_20829);
  nand g46732 (n_16497, n_17748, n_16496);
  nand g46733 (n_16334, n_17749, n_16333);
  nand g46734 (n_20814, \data_stack_mem[2] [3], n_16402);
  nand g46735 (n_20820, \data_stack_mem[3] [2], n_16322);
  nand g46736 (n_24507, n_16221, n_16228);
  or g46737 (n_24508, n_16221, n_16228);
  nand g46738 (n_16229, n_24507, n_24508);
  nand g46739 (n_16656, n_17738, n_16655);
  nand g46740 (n_17424, n_18486, n_18487);
  nand g46741 (n_20920, n_20918, n_20919);
  or g46742 (n_20808, \data_stack_mem[2] [3], wc302);
  not gc302 (wc302, n_16377);
  nand g46743 (n_24509, n_16244, n_16253);
  or g46744 (n_24510, n_16244, n_16253);
  nand g46745 (n_16254, n_24509, n_24510);
  or g46746 (n_17700, n_20848, n_16178);
  or g46749 (n_19448, n_16681, n_16731);
  or g46750 (n_22999, wc303, n_16683);
  not gc303 (wc303, n_17294);
  or g46752 (n_19435, n_16683, n_16680);
  nand g46753 (n_19129, n_19127, n_19128);
  nand g46754 (n_16419, n_17760, n_16418);
  or g46756 (n_20937, \data_stack_mem[8] [1], wc304);
  not gc304 (wc304, n_16214);
  nand g46757 (n_19117, n_19115, n_19116);
  nand g46758 (n_23047, n_16228, n_17348);
  nand g46759 (n_24511, n_16292, n_16294);
  or g46760 (n_24512, n_16292, n_16294);
  nand g46761 (n_16295, n_24511, n_24512);
  nand g46762 (n_23062, n_16253, n_17409);
  nand g46763 (n_16297, n_19590, n_23041);
  nand g46764 (n_16315, n_20712, n_23050);
  or g46765 (n_20758, n_16296, wc305);
  not gc305 (wc305, n_16322);
  or g46766 (n_20757, n_16268, n_16322);
  nand g46767 (n_24513, n_16318, n_16320);
  or g46768 (n_24514, n_16318, n_16320);
  nand g46769 (n_16321, n_24513, n_24514);
  nand g46770 (n_23041, n_17450, n_16227);
  nand g46771 (n_16377, n_20718, n_23053);
  or g46772 (n_17695, n_20782, n_16178);
  nand g46773 (n_20848, n_20846, n_20847);
  nand g46774 (n_17027, n_19566, n_19567);
  nand g46775 (n_16953, n_19155, n_19156);
  or g46776 (n_17131, n_19926, n_19927);
  nand g46777 (n_16261, n_17739, n_16260);
  nand g46778 (n_24515, n_16246, n_16252);
  or g46779 (n_24516, n_16246, n_16252);
  nand g46780 (n_16253, n_24515, n_24516);
  or g46781 (n_16184, n_16183, wc306);
  not gc306 (wc306, n_18226);
  or g46782 (n_17146, n_20502, n_20503);
  nand g46783 (n_17028, n_19572, n_19573);
  or g46784 (n_17126, n_19686, n_19687);
  nand g46786 (n_17029, n_19578, n_19579);
  nand g46787 (n_17011, n_19482, n_19483);
  nand g46788 (n_16954, n_19161, n_19162);
  or g46790 (n_20828, \data_stack_mem[7] [1], wc307);
  not gc307 (wc307, n_16240);
  or g46791 (n_20919, wc308, n_16542);
  not gc308 (wc308, n_17310);
  or g46792 (n_20918, n_17310, wc309);
  not gc309 (wc309, n_16542);
  or g46793 (n_17147, n_20550, n_20551);
  nand g46794 (n_16955, n_19167, n_19168);
  nand g46795 (n_17012, n_19488, n_19489);
  or g46796 (n_20838, n_16210, wc310);
  not gc310 (wc310, n_16232);
  or g46797 (n_20829, wc311, n_16240);
  not gc311 (wc311, \data_stack_mem[7] [1]);
  nand g46798 (n_17030, n_19584, n_19585);
  or g46799 (n_20839, \data_stack_mem[7] [1], n_20837);
  or g46800 (n_17749, n_19042, n_16179);
  nand g46801 (n_16999, n_19317, n_19318);
  nand g46802 (n_16956, n_19173, n_19174);
  nand g46804 (n_16402, n_20724, n_23056);
  nand g46805 (n_17013, n_19494, n_19495);
  nand g46806 (n_24517, n_16147, n_16170);
  or g46807 (n_24518, n_16147, n_16170);
  nand g46808 (n_16171, n_24517, n_24518);
  nand g46809 (n_16957, n_19179, n_19180);
  nand g46810 (n_17000, n_19323, n_19324);
  nand g46811 (n_16958, n_19185, n_19186);
  nand g46812 (n_20803, n_17328, n_20802);
  or g46813 (n_17128, n_19782, n_19783);
  nand g46814 (n_17001, n_19329, n_19330);
  nand g46815 (n_16959, n_19191, n_19192);
  nand g46816 (n_17014, n_19500, n_19501);
  nand g46818 (n_16960, n_19197, n_19198);
  nand g46819 (n_17002, n_19335, n_19336);
  or g46820 (n_20910, \data_stack_mem[7] [1], wc312);
  not gc312 (wc312, n_16232);
  nand g46821 (n_17015, n_19506, n_19507);
  nand g46822 (n_16961, n_19203, n_19204);
  nand g46823 (n_17003, n_19341, n_19342);
  nand g46824 (n_16322, n_19596, n_23044);
  nand g46825 (n_16964, n_19209, n_19210);
  nand g46826 (n_20857, n_20855, n_20856);
  or g46827 (n_17136, n_20118, n_20119);
  nand g46828 (n_17004, n_19347, n_19348);
  nand g46829 (n_16965, n_19215, n_19216);
  nand g46830 (n_17016, n_19512, n_19513);
  nand g46831 (n_20797, n_17397, n_20796);
  or g46832 (n_17140, n_20646, n_20647);
  nand g46833 (n_16966, n_19221, n_19222);
  nand g46834 (n_17005, n_19353, n_19354);
  or g46835 (n_17144, n_20406, n_20407);
  or g46836 (n_16788, n_16183, wc313);
  not gc313 (wc313, n_18085);
  nand g46837 (n_16967, n_19227, n_19228);
  or g46838 (n_16418, n_16183, wc314);
  not gc314 (wc314, n_18247);
  or g46839 (n_16244, n_20752, wc315);
  not gc315 (wc315, n_16154);
  or g46840 (n_17748, n_19012, n_16179);
  nand g46841 (n_17006, n_19359, n_19360);
  nand g46842 (n_16968, n_19233, n_19234);
  nand g46843 (n_17017, n_19518, n_19519);
  or g46844 (n_17750, n_19072, n_16179);
  or g46845 (n_17130, n_19878, n_19879);
  nand g46846 (n_16969, n_19239, n_19240);
  or g46847 (n_17760, n_19102, n_16179);
  nand g46848 (n_17007, n_19365, n_19366);
  or g46849 (n_17135, n_20598, n_20599);
  nand g46850 (n_16970, n_19245, n_19246);
  or g46851 (n_17738, n_18949, n_16179);
  nand g46852 (n_17018, n_19524, n_19525);
  nand g46854 (n_16971, n_19251, n_19252);
  or g46855 (n_17145, n_20454, n_20455);
  nand g46856 (n_17019, n_19530, n_19531);
  or g46857 (n_16219, n_20746, wc316);
  not gc316 (wc316, n_16154);
  or g46858 (n_17705, n_20791, n_16178);
  nand g46859 (n_16972, n_19257, n_19258);
  or g46860 (n_17133, n_20022, n_20023);
  nand g46862 (n_17022, n_19536, n_19537);
  nand g46863 (n_24519, n_16223, n_16227);
  or g46864 (n_24520, n_16223, n_16227);
  nand g46865 (n_16228, n_24519, n_24520);
  or g46866 (n_17134, n_20070, n_20071);
  or g46867 (n_17141, n_20694, n_20695);
  or g46868 (n_17127, n_19734, n_19735);
  or g46869 (n_17142, n_20310, n_20311);
  nand g46870 (n_17023, n_19542, n_19543);
  or g46871 (n_17129, n_19830, n_19831);
  nand g46872 (n_16683, n_17908, n_22996);
  or g46873 (n_17139, n_20262, n_20263);
  or g46874 (n_17143, n_20358, n_20359);
  nand g46875 (n_17024, n_19548, n_19549);
  or g46876 (n_17132, n_19974, n_19975);
  nand g46877 (n_16731, n_18106, n_23005);
  or g46878 (n_17138, n_20214, n_20215);
  nand g46879 (n_17025, n_19554, n_19555);
  nand g46880 (n_23050, n_16252, n_17415);
  or g46881 (n_17137, n_20166, n_20167);
  nand g46882 (n_17026, n_19560, n_19561);
  or g46883 (n_17668, n_20773, n_16178);
  nand g46884 (n_19360, \data_stack_mem[9] [2], n_16998);
  nand g46885 (n_19366, data_parity_mem[9], n_16998);
  nand g46886 (n_20725, n_17378, n_20724);
  nand g46887 (n_17033, n_19371, n_19372);
  nand g46888 (n_19354, \data_stack_mem[9] [6], n_16998);
  or g46889 (n_21014, n_16484, n_16458);
  nand g46890 (n_19348, \data_stack_mem[9] [0], n_16998);
  nand g46891 (n_19342, \data_stack_mem[9] [4], n_16998);
  nand g46892 (n_17034, n_19377, n_19378);
  nand g46893 (n_23044, n_17429, n_16251);
  nand g46894 (n_19336, \data_stack_mem[9] [7], n_16998);
  nand g46895 (n_19330, \data_stack_mem[9] [5], n_16998);
  nand g46896 (n_17035, n_19383, n_19384);
  nand g46897 (n_19324, \data_stack_mem[9] [1], n_16998);
  nand g46898 (n_19318, \data_stack_mem[9] [3], n_16998);
  or g46899 (n_20263, n_20260, n_20261);
  nand g46900 (n_16996, n_19311, n_19312);
  nand g46901 (n_16995, n_19305, n_19306);
  nand g46902 (n_16994, n_19299, n_19300);
  nand g46903 (n_17036, n_19389, n_19390);
  nand g46904 (n_16993, n_19293, n_19294);
  nand g46905 (n_16992, n_19287, n_19288);
  nand g46906 (n_17037, n_19395, n_19396);
  or g46907 (n_20215, n_20212, n_20213);
  or g46908 (n_20359, n_20356, n_20357);
  nand g46909 (n_23005, n_17427, n_16617);
  nand g46910 (n_16991, n_19281, n_19282);
  nand g46911 (n_17038, n_19401, n_19402);
  nand g46912 (n_16990, n_19275, n_19276);
  nand g46913 (n_16989, n_19269, n_19270);
  nand g46914 (n_16988, n_19263, n_19264);
  nand g46915 (n_19258, data_parity_mem[3], n_16963);
  nand g46916 (n_19252, \data_stack_mem[3] [2], n_16963);
  nand g46917 (n_19246, \data_stack_mem[3] [0], n_16963);
  nand g46918 (n_17039, n_19407, n_19408);
  nand g46919 (n_24521, n_16149, n_16169);
  or g46920 (n_20837, n_16149, n_16169);
  nand g46921 (n_16170, n_24521, n_20837);
  or g46922 (n_20932, \data_stack_mem[2] [4], wc317);
  not gc317 (wc317, n_16484);
  nand g46923 (n_19240, \data_stack_mem[3] [4], n_16963);
  nand g46924 (n_19234, \data_stack_mem[3] [5], n_16963);
  nand g46925 (n_19228, \data_stack_mem[3] [6], n_16963);
  nand g46926 (n_17040, n_19413, n_19414);
  nand g46927 (n_19222, \data_stack_mem[3] [7], n_16963);
  nand g46928 (n_19216, \data_stack_mem[3] [1], n_16963);
  nand g46929 (n_19210, \data_stack_mem[3] [3], n_16963);
  nand g46930 (n_17041, n_19419, n_19420);
  nand g46931 (n_19204, data_parity_mem[1], n_16952);
  nand g46932 (n_19198, \data_stack_mem[1] [7], n_16952);
  nand g46933 (n_19192, \data_stack_mem[1] [0], n_16952);
  nand g46934 (n_19186, \data_stack_mem[1] [6], n_16952);
  nand g46935 (n_19180, \data_stack_mem[1] [4], n_16952);
  nand g46936 (n_19483, \data_stack_mem[7] [2], n_17010);
  nand g46937 (n_19174, \data_stack_mem[1] [3], n_16952);
  nand g46938 (n_19489, \data_stack_mem[7] [0], n_17010);
  nand g46939 (n_19168, \data_stack_mem[1] [1], n_16952);
  nand g46940 (n_19495, \data_stack_mem[7] [7], n_17010);
  or g46942 (n_20407, n_20404, n_20405);
  or g46943 (n_20796, \data_stack_mem[6] [1], wc318);
  not gc318 (wc318, n_16216);
  or g46944 (n_20167, n_20164, n_20165);
  nand g46945 (n_19162, \data_stack_mem[1] [2], n_16952);
  nand g46946 (n_19501, \data_stack_mem[7] [5], n_17010);
  nand g46947 (n_19507, data_parity_mem[7], n_17010);
  nand g46948 (n_19513, \data_stack_mem[7] [4], n_17010);
  nand g46949 (n_19519, \data_stack_mem[7] [3], n_17010);
  nand g46950 (n_19156, \data_stack_mem[1] [5], n_16952);
  nand g46952 (n_19525, \data_stack_mem[7] [1], n_17010);
  nand g46953 (n_19531, \data_stack_mem[7] [6], n_17010);
  nand g46954 (n_19537, \data_stack_mem[5] [0], n_17021);
  nand g46955 (n_19543, \data_stack_mem[5] [1], n_17021);
  nand g46956 (n_22996, n_17443, n_16643);
  or g46957 (n_20071, n_20068, n_20069);
  nand g46958 (n_19555, \data_stack_mem[5] [3], n_17021);
  or g46959 (n_19102, wc319, n_19101);
  not gc319 (wc319, n_16391);
  or g46960 (n_20455, n_20452, n_20453);
  nand g46961 (n_19561, \data_stack_mem[5] [5], n_17021);
  nand g46962 (n_19567, \data_stack_mem[5] [6], n_17021);
  nand g46963 (n_19573, \data_stack_mem[5] [7], n_17021);
  nand g46964 (n_19579, data_parity_mem[5], n_17021);
  nand g46965 (n_19585, \data_stack_mem[5] [4], n_17021);
  or g46966 (n_17080, n_19638, n_19639);
  or g46967 (n_20503, n_20500, n_20501);
  nand g46968 (n_20746, n_17405, n_20745);
  or g46969 (n_19687, n_19684, n_19685);
  or g46971 (n_19126, n_16643, n_16594);
  or g46972 (n_19735, n_19732, n_19733);
  or g46973 (n_20551, n_20548, n_20549);
  or g46974 (n_19783, n_19780, n_19781);
  nand g46975 (n_20791, n_20789, n_20790);
  nand g46976 (n_16915, n_18729, n_18730);
  nand g46977 (n_20719, n_17365, n_20718);
  nand g46978 (n_16914, n_18723, n_18724);
  nand g46979 (n_16913, n_18717, n_18718);
  nand g46980 (n_24523, n_16248, n_16251);
  or g46981 (n_24524, n_16248, n_16251);
  nand g46982 (n_16252, n_24523, n_24524);
  nand g46983 (n_16912, n_18711, n_18712);
  nand g46984 (n_16911, n_18705, n_18706);
  nand g46985 (n_16910, n_18699, n_18700);
  nand g46986 (n_16909, n_18693, n_18694);
  or g46987 (n_19831, n_19828, n_19829);
  or g46988 (n_20599, n_20596, n_20597);
  or g46990 (n_19115, n_16595, n_16617);
  or g46991 (n_19042, wc320, n_19041);
  not gc320 (wc320, n_16306);
  or g46992 (n_16333, n_16183, wc321);
  not gc321 (wc321, n_18202);
  nand g46993 (n_16908, n_18687, n_18688);
  or g46994 (n_20119, n_20116, n_20117);
  nand g46995 (n_20782, n_20780, n_20781);
  or g46996 (n_19879, n_19876, n_19877);
  or g46997 (n_16246, n_20713, wc322);
  not gc322 (wc322, n_16156);
  or g46998 (n_20847, wc323, n_16369);
  not gc323 (wc323, n_16351);
  or g46999 (n_20846, n_16351, wc324);
  not gc324 (wc324, n_16369);
  or g47000 (n_19012, wc325, n_19011);
  not gc325 (wc325, n_16471);
  nand g47001 (n_20752, n_17409, n_20751);
  nand g47002 (n_23053, n_17365, n_16294);
  or g47003 (n_16496, n_16183, wc326);
  not gc326 (wc326, n_18181);
  or g47004 (n_20647, n_20644, n_20645);
  or g47005 (n_19927, n_19924, n_19925);
  or g47006 (n_20802, wc327, n_16241);
  not gc327 (wc327, \data_stack_mem[6] [1]);
  or g47008 (n_17646, n_20734, n_16178);
  or g47009 (n_19975, n_19972, n_19973);
  or g47010 (n_20311, n_20308, n_20309);
  nand g47011 (n_24525, n_17461, n_16541);
  or g47012 (n_24526, n_17461, n_16541);
  nand g47013 (n_16542, n_24525, n_24526);
  or g47014 (n_20695, n_20692, n_20693);
  or g47015 (n_16221, n_20707, wc328);
  not gc328 (wc328, n_16156);
  or g47016 (n_19072, wc329, n_19071);
  not gc329 (wc329, n_16785);
  or g47018 (n_20855, n_16195, wc330);
  not gc330 (wc330, n_16213);
  or g47019 (n_20856, wc331, n_16213);
  not gc331 (wc331, n_16195);
  or g47020 (n_20023, n_20020, n_20021);
  nand g47021 (n_23056, n_17378, n_16320);
  nand g47023 (n_17751, n_18159, n_18160);
  nand g47024 (n_23035, n_23033, n_23034);
  or g47025 (n_17739, n_18982, n_16179);
  or g47026 (n_16260, n_16183, wc332);
  not gc332 (wc332, n_18148);
  nand g47027 (n_20773, n_20771, n_20772);
  or g47028 (n_16227, wc333, n_19465);
  not gc333 (wc333, n_19464);
  or g47029 (n_18949, wc334, n_18948);
  not gc334 (wc334, n_16628);
  or g47030 (n_16655, n_16183, wc335);
  not gc335 (wc335, n_18127);
  nand g47031 (n_18486, n_16183, n_17752);
  nand g47032 (n_19549, \data_stack_mem[5] [2], n_17021);
  nand g47034 (n_20734, n_20732, n_20733);
  or g47035 (n_19686, n_19682, n_19683);
  or g47036 (n_20070, n_20066, n_20067);
  nand g47040 (n_24527, n_16153, n_16168);
  or g47041 (n_24528, n_16153, n_16168);
  nand g47042 (n_16169, n_24527, n_24528);
  nand g47043 (n_16120, n_18609, n_18610);
  nand g47044 (n_19396, \data_stack_mem[4] [0], n_17032);
  or g47048 (n_19974, n_19970, n_19971);
  or g47049 (n_20166, n_20162, n_20163);
  nand g47051 (n_19464, n_17654, n_16225);
  or g47053 (n_17757, n_18523, n_16179);
  or g47054 (n_19830, n_19826, n_19827);
  nand g47055 (n_16251, n_20700, n_20701);
  or g47056 (n_17752, wc336, n_16500);
  not gc336 (wc336, n_18160);
  or g47058 (n_20502, n_20498, n_20499);
  nand g47060 (n_18541, n_18538, n_18539);
  nand g47062 (n_19294, \data_stack_mem[6] [0], n_16987);
  or g47063 (n_20406, n_20402, n_20403);
  nand g47066 (n_19264, \data_stack_mem[6] [5], n_16987);
  or g47067 (n_19926, n_19922, n_19923);
  nand g47068 (n_16123, n_18615, n_18616);
  nand g47070 (n_19390, data_parity_mem[4], n_17032);
  or g47071 (n_20745, \data_stack_mem[5] [1], wc337);
  not gc337 (wc337, n_16218);
  nand g47072 (n_16126, n_18621, n_18622);
  or g47073 (n_19639, n_19636, n_19637);
  or g47074 (n_20751, wc338, n_16243);
  not gc338 (wc338, \data_stack_mem[5] [1]);
  or g47075 (n_20790, wc339, n_16282);
  not gc339 (wc339, n_16264);
  or g47076 (n_20646, n_20642, n_20643);
  or g47077 (n_20789, n_16264, wc340);
  not gc340 (wc340, n_16282);
  nand g47078 (n_16129, n_18627, n_18628);
  nand g47079 (n_16916, n_18735, n_18736);
  or g47080 (n_19638, n_19634, n_19635);
  nand g47081 (n_16132, n_18633, n_18634);
  or g47084 (n_17021, n_17009, wc341);
  not gc341 (wc341, n_19477);
  nand g47087 (n_16917, n_18741, n_18742);
  or g47089 (n_20118, n_20114, n_20115);
  nand g47090 (n_19270, \data_stack_mem[6] [4], n_16987);
  or g47091 (n_20772, wc342, n_16604);
  not gc342 (wc342, n_16586);
  or g47092 (n_20771, n_16586, wc343);
  not gc343 (wc343, n_16604);
  nand g47094 (n_16918, n_18747, n_18748);
  nand g47095 (n_19300, \data_stack_mem[6] [1], n_16987);
  nand g47096 (n_19372, \data_stack_mem[4] [5], n_17032);
  nand g47098 (n_16919, n_18753, n_18754);
  or g47100 (n_17010, n_17009, wc344);
  not gc344 (wc344, n_19474);
  nand g47102 (n_16920, n_18759, n_18760);
  nand g47103 (n_20713, n_17415, n_20712);
  nand g47104 (n_19276, \data_stack_mem[6] [3], n_16987);
  nand g47106 (n_16921, n_18765, n_18766);
  nand g47107 (n_19384, \data_stack_mem[4] [7], n_17032);
  or g47109 (n_18159, n_16145, wc345);
  not gc345 (wc345, n_16500);
  nand g47110 (n_16922, n_18771, n_18772);
  nand g47111 (n_16899, n_18639, n_18640);
  or g47112 (n_20454, n_20450, n_20451);
  nand g47114 (n_16900, n_18645, n_18646);
  or g47115 (n_19878, n_19874, n_19875);
  nand g47116 (n_16923, n_18777, n_18778);
  nand g47117 (n_16901, n_18651, n_18652);
  nand g47118 (n_19306, \data_stack_mem[6] [6], n_16987);
  or g47119 (n_20022, n_20018, n_20019);
  nand g47120 (n_16902, n_18657, n_18658);
  nand g47122 (n_19420, \data_stack_mem[4] [4], n_17032);
  nand g47124 (n_16903, n_18663, n_18664);
  nand g47127 (n_16213, n_24529, n_24530);
  or g47128 (n_19782, n_19778, n_19779);
  nand g47129 (n_16904, n_18669, n_18670);
  nand g47132 (n_16905, n_18675, n_18676);
  nand g47133 (n_19282, \data_stack_mem[6] [2], n_16987);
  nand g47135 (n_19378, \data_stack_mem[4] [6], n_17032);
  or g47136 (n_20781, wc346, n_16447);
  not gc346 (wc346, n_16429);
  or g47137 (n_20780, n_16429, wc347);
  not gc347 (wc347, n_16447);
  nand g47138 (n_16906, n_18681, n_18682);
  or g47141 (n_20550, n_20546, n_20547);
  nand g47145 (n_19402, \data_stack_mem[4] [2], n_17032);
  nand g47147 (n_19414, \data_stack_mem[4] [1], n_17032);
  nand g47150 (n_16369, n_24531, n_24532);
  or g47151 (n_20262, n_20258, n_20259);
  or g47152 (n_16998, n_19144, n_16951);
  nand g47156 (n_16617, n_18546, n_18547);
  or g47157 (n_20310, n_20306, n_20307);
  nand g47159 (n_24533, n_16505, n_16540);
  or g47160 (n_24534, n_16505, n_16540);
  nand g47161 (n_16541, n_24533, n_24534);
  or g47163 (n_19734, n_19730, n_19731);
  or g47165 (n_20358, n_20354, n_20355);
  or g47167 (n_20718, \data_stack_mem[2] [2], wc348);
  not gc348 (wc348, n_16291);
  or g47168 (n_20598, n_20594, n_20595);
  or g47169 (n_20694, n_20690, n_20691);
  or g47172 (n_20214, n_20210, n_20211);
  nand g47174 (n_19288, data_parity_mem[6], n_16987);
  nand g47175 (n_20707, n_17348, n_20706);
  nand g47177 (n_19408, \data_stack_mem[4] [3], n_17032);
  nand g47179 (n_16111, n_18591, n_18592);
  nand g47180 (n_16643, n_17905, n_22993);
  nand g47181 (n_19312, \data_stack_mem[6] [7], n_16987);
  nand g47182 (n_16114, n_18597, n_18598);
  nand g47184 (n_20724, \data_stack_mem[2] [2], n_16317);
  nand g47185 (n_16117, n_18603, n_18604);
  nand g47186 (n_16317, n_19425, n_23038);
  or g47187 (n_22573, wc349, n_16124);
  not gc349 (wc349, \out_fifo[2][1] [7]);
  or g47188 (n_22570, wc350, n_16124);
  not gc350 (wc350, \out_fifo[2][1] [5]);
  nand g47189 (n_19591, n_17450, n_19590);
  or g47190 (n_22567, wc351, n_16124);
  not gc351 (wc351, \out_fifo[2][1] [8]);
  or g47191 (n_22564, wc352, n_16124);
  not gc352 (wc352, \out_fifo[2][1] [6]);
  or g47192 (n_22561, wc353, n_16130);
  not gc353 (wc353, \out_fifo[1][1] [8]);
  or g47193 (n_22558, wc354, n_16130);
  not gc354 (wc354, \out_fifo[1][1] [7]);
  or g47194 (n_22555, wc355, n_16130);
  not gc355 (wc355, \out_fifo[1][1] [6]);
  or g47196 (n_22552, wc356, n_16130);
  not gc356 (wc356, \out_fifo[1][1] [5]);
  or g47197 (n_22549, wc357, n_16109);
  not gc357 (wc357, \out_fifo[7][1] [6]);
  or g47198 (n_22546, wc358, n_16109);
  not gc358 (wc358, \out_fifo[7][1] [7]);
  or g47199 (n_22543, wc359, n_16109);
  not gc359 (wc359, \out_fifo[7][1] [5]);
  or g47200 (n_22540, wc360, n_16109);
  not gc360 (wc360, \out_fifo[7][1] [8]);
  nand g47201 (n_20068, n_20062, n_20063);
  or g47202 (n_22528, wc361, n_16130);
  not gc361 (wc361, \out_fifo[1][0] [8]);
  or g47203 (n_22522, wc362, n_16127);
  not gc362 (wc362, \out_fifo[4][0] [8]);
  nand g47205 (n_20067, n_20060, n_20061);
  or g47206 (n_22516, wc363, n_16124);
  not gc363 (wc363, \out_fifo[2][0] [8]);
  or g47207 (n_22510, wc364, n_16121);
  not gc364 (wc364, \out_fifo[0][0] [8]);
  or g47208 (n_22504, wc365, n_16118);
  not gc365 (wc365, \out_fifo[6][0] [8]);
  or g47209 (n_22498, wc366, n_16115);
  not gc366 (wc366, \out_fifo[3][0] [8]);
  nand g47210 (n_20066, n_20058, n_20059);
  nand g47211 (n_20305, n_20296, n_20297);
  or g47212 (n_18947, n_18945, n_18946);
  nand g47213 (n_20065, n_20056, n_20057);
  or g47214 (n_22492, wc367, n_16112);
  not gc367 (wc367, \out_fifo[5][0] [8]);
  or g47215 (n_22486, wc368, n_16109);
  not gc368 (wc368, \out_fifo[7][0] [8]);
  or g47216 (n_22399, wc369, n_16130);
  not gc369 (wc369, \out_fifo[1][0] [7]);
  or g47217 (n_22393, wc370, n_16127);
  not gc370 (wc370, \out_fifo[4][0] [7]);
  nand g47218 (n_20306, n_20298, n_20299);
  nand g47219 (n_19465, n_19462, n_19463);
  or g47220 (n_22576, wc371, n_16121);
  not gc371 (wc371, \out_fifo[0][1] [6]);
  or g47221 (n_22387, wc372, n_16124);
  not gc372 (wc372, \out_fifo[2][0] [7]);
  or g47222 (n_22381, wc373, n_16121);
  not gc373 (wc373, \out_fifo[0][0] [7]);
  or g47223 (n_22375, wc374, n_16118);
  not gc374 (wc374, \out_fifo[6][0] [7]);
  or g47224 (n_22369, wc375, n_16115);
  not gc375 (wc375, \out_fifo[3][0] [7]);
  or g47225 (n_22363, wc376, n_16112);
  not gc376 (wc376, \out_fifo[5][0] [7]);
  or g47226 (n_22357, wc377, n_16109);
  not gc377 (wc377, \out_fifo[7][0] [7]);
  or g47227 (n_22333, wc378, n_16130);
  not gc378 (wc378, \out_fifo[1][0] [6]);
  or g47228 (n_22327, wc379, n_16127);
  not gc379 (wc379, \out_fifo[4][0] [6]);
  or g47229 (n_22321, wc380, n_16124);
  not gc380 (wc380, \out_fifo[2][0] [6]);
  or g47230 (n_22315, wc381, n_16121);
  not gc381 (wc381, \out_fifo[0][0] [6]);
  nand g47231 (n_16291, n_19470, n_19471);
  or g47232 (n_22309, wc382, n_16118);
  not gc382 (wc382, \out_fifo[6][0] [6]);
  or g47233 (n_22303, wc383, n_16115);
  not gc383 (wc383, \out_fifo[3][0] [6]);
  nand g47234 (n_20307, n_20300, n_20301);
  or g47235 (n_22297, wc384, n_16112);
  not gc384 (wc384, \out_fifo[5][0] [6]);
  or g47236 (n_22291, wc385, n_16109);
  not gc385 (wc385, \out_fifo[7][0] [6]);
  or g47237 (n_22579, wc386, n_16121);
  not gc386 (wc386, \out_fifo[0][1] [7]);
  or g47239 (n_22177, wc387, n_16130);
  not gc387 (wc387, \out_fifo[1][0] [5]);
  or g47240 (n_22171, wc388, n_16127);
  not gc388 (wc388, \out_fifo[4][0] [5]);
  or g47241 (n_22582, wc389, n_16121);
  not gc389 (wc389, \out_fifo[0][1] [8]);
  or g47243 (n_22165, wc390, n_16124);
  not gc390 (wc390, \out_fifo[2][0] [5]);
  or g47244 (n_22159, wc391, n_16121);
  not gc391 (wc391, \out_fifo[0][0] [5]);
  or g47245 (n_22153, wc392, n_16118);
  not gc392 (wc392, \out_fifo[6][0] [5]);
  or g47247 (n_22585, wc393, n_16121);
  not gc393 (wc393, \out_fifo[0][1] [5]);
  nand g47248 (n_20113, n_20104, n_20105);
  or g47249 (n_18981, n_18979, n_18980);
  or g47251 (n_22147, wc394, n_16115);
  not gc394 (wc394, \out_fifo[3][0] [5]);
  or g47252 (n_22141, wc395, n_16112);
  not gc395 (wc395, \out_fifo[5][0] [5]);
  or g47253 (n_22588, wc396, n_16115);
  not gc396 (wc396, \out_fifo[3][1] [7]);
  or g47254 (n_22135, wc397, n_16109);
  not gc397 (wc397, \out_fifo[7][0] [5]);
  or g47255 (n_21919, wc398, n_16130);
  not gc398 (wc398, \out_fifo[1][0] [4]);
  or g47256 (n_21913, wc399, n_16127);
  not gc399 (wc399, \out_fifo[4][0] [4]);
  or g47257 (n_21907, wc400, n_16124);
  not gc400 (wc400, \out_fifo[2][0] [4]);
  or g47258 (n_22591, wc401, n_16115);
  not gc401 (wc401, \out_fifo[3][1] [6]);
  or g47259 (n_21901, wc402, n_16121);
  not gc402 (wc402, \out_fifo[0][0] [4]);
  or g47260 (n_21895, wc403, n_16118);
  not gc403 (wc403, \out_fifo[6][0] [4]);
  or g47261 (n_21889, wc404, n_16115);
  not gc404 (wc404, \out_fifo[3][0] [4]);
  or g47262 (n_21883, wc405, n_16112);
  not gc405 (wc405, \out_fifo[5][0] [4]);
  nand g47263 (n_20020, n_20014, n_20015);
  or g47264 (n_21877, wc406, n_16109);
  not gc406 (wc406, \out_fifo[7][0] [4]);
  or g47265 (n_21721, wc407, n_16130);
  not gc407 (wc407, \out_fifo[1][0] [3]);
  nand g47266 (n_20019, n_20012, n_20013);
  or g47267 (n_21715, wc408, n_16127);
  not gc408 (wc408, \out_fifo[4][0] [3]);
  or g47268 (n_21709, wc409, n_16124);
  not gc409 (wc409, \out_fifo[2][0] [3]);
  or g47269 (n_21703, wc410, n_16121);
  not gc410 (wc410, \out_fifo[0][0] [3]);
  or g47270 (n_21697, wc411, n_16118);
  not gc411 (wc411, \out_fifo[6][0] [3]);
  or g47271 (n_21691, wc412, n_16115);
  not gc412 (wc412, \out_fifo[3][0] [3]);
  nand g47272 (n_20018, n_20010, n_20011);
  or g47273 (n_21685, wc413, n_16112);
  not gc413 (wc413, \out_fifo[5][0] [3]);
  or g47274 (n_22594, wc414, n_16115);
  not gc414 (wc414, \out_fifo[3][1] [5]);
  nand g47275 (n_17125, n_16116, n_18103);
  or g47276 (n_21679, wc415, n_16109);
  not gc415 (wc415, \out_fifo[7][0] [3]);
  or g47277 (n_21424, wc416, n_16130);
  not gc416 (wc416, \out_fifo[1][0] [2]);
  nand g47278 (n_20308, n_20302, n_20303);
  or g47279 (n_21418, wc417, n_16127);
  not gc417 (wc417, \out_fifo[4][0] [2]);
  or g47280 (n_21412, wc418, n_16124);
  not gc418 (wc418, \out_fifo[2][0] [2]);
  or g47281 (n_21406, wc419, n_16121);
  not gc419 (wc419, \out_fifo[0][0] [2]);
  or g47282 (n_22597, wc420, n_16115);
  not gc420 (wc420, \out_fifo[3][1] [8]);
  nand g47284 (n_20017, n_20008, n_20009);
  or g47285 (n_21400, wc421, n_16118);
  not gc421 (wc421, \out_fifo[6][0] [2]);
  or g47286 (n_21394, wc422, n_16115);
  not gc422 (wc422, \out_fifo[3][0] [2]);
  or g47287 (n_21388, wc423, n_16112);
  not gc423 (wc423, \out_fifo[5][0] [2]);
  nand g47288 (n_20114, n_20106, n_20107);
  or g47289 (n_19070, n_19068, n_19069);
  or g47290 (n_21382, wc424, n_16109);
  not gc424 (wc424, \out_fifo[7][0] [2]);
  or g47291 (n_21160, wc425, n_16130);
  not gc425 (wc425, \out_fifo[1][0] [1]);
  or g47292 (n_21154, wc426, n_16127);
  not gc426 (wc426, \out_fifo[4][0] [1]);
  or g47293 (n_21148, wc427, n_16124);
  not gc427 (wc427, \out_fifo[2][0] [1]);
  or g47294 (n_21142, wc428, n_16121);
  not gc428 (wc428, \out_fifo[0][0] [1]);
  or g47295 (n_21136, wc429, n_16118);
  not gc429 (wc429, \out_fifo[6][0] [1]);
  or g47296 (n_21130, wc430, n_16115);
  not gc430 (wc430, \out_fifo[3][0] [1]);
  or g47297 (n_21124, wc431, n_16112);
  not gc431 (wc431, \out_fifo[5][0] [1]);
  or g47298 (n_21118, wc432, n_16109);
  not gc432 (wc432, \out_fifo[7][0] [1]);
  or g47299 (n_22600, wc433, n_16112);
  not gc433 (wc433, \out_fifo[5][1] [6]);
  nand g47300 (n_20692, n_20686, n_20687);
  nand g47301 (n_20691, n_20684, n_20685);
  nand g47302 (n_20690, n_20682, n_20683);
  nand g47303 (n_20689, n_20680, n_20681);
  nand g47304 (n_20115, n_20108, n_20109);
  or g47306 (n_18592, wc434, n_16109);
  not gc434 (wc434, \out_fifo[7][2] [6]);
  or g47308 (n_18598, wc435, n_16112);
  not gc435 (wc435, \out_fifo[5][2] [6]);
  or g47309 (n_18603, wc436, n_16116);
  not gc436 (wc436, n_16108);
  or g47310 (n_18604, wc437, n_16115);
  not gc437 (wc437, \out_fifo[3][2] [6]);
  or g47311 (n_22603, wc438, n_16112);
  not gc438 (wc438, \out_fifo[5][1] [7]);
  or g47312 (n_20733, wc439, n_16784);
  not gc439 (wc439, n_16771);
  or g47313 (n_20732, n_16771, wc440);
  not gc440 (wc440, n_16784);
  or g47315 (n_18610, wc441, n_16118);
  not gc441 (wc441, \out_fifo[6][2] [6]);
  nand g47316 (n_20116, n_20110, n_20111);
  nand g47320 (n_16604, n_24535, n_24536);
  nand g47321 (n_19972, n_19966, n_19967);
  or g47322 (n_22606, wc442, n_16112);
  not gc442 (wc442, \out_fifo[5][1] [8]);
  or g47323 (n_18523, n_18521, n_18522);
  nand g47326 (n_16447, n_24537, n_24538);
  or g47328 (n_18616, wc443, n_16121);
  not gc443 (wc443, \out_fifo[0][2] [6]);
  nand g47329 (n_19971, n_19964, n_19965);
  or g47330 (n_22609, wc444, n_16112);
  not gc444 (wc444, \out_fifo[5][1] [5]);
  nand g47331 (n_19970, n_19962, n_19963);
  nand g47332 (n_19969, n_19960, n_19961);
  or g47333 (n_22612, wc445, n_16118);
  not gc445 (wc445, \out_fifo[6][1] [7]);
  or g47334 (n_22615, wc446, n_16118);
  not gc446 (wc446, \out_fifo[6][1] [5]);
  or g47336 (n_18622, wc447, n_16124);
  not gc447 (wc447, \out_fifo[2][2] [6]);
  or g47338 (n_22618, wc448, n_16118);
  not gc448 (wc448, \out_fifo[6][1] [6]);
  or g47339 (n_18628, wc449, n_16127);
  not gc449 (wc449, \out_fifo[4][2] [6]);
  or g47341 (n_18634, wc450, n_16130);
  not gc450 (wc450, \out_fifo[1][2] [6]);
  nand g47343 (n_20644, n_20638, n_20639);
  nand g47344 (n_20643, n_20636, n_20637);
  or g47345 (n_22621, wc451, n_16118);
  not gc451 (wc451, \out_fifo[6][1] [8]);
  or g47346 (n_19010, n_19008, n_19009);
  nand g47347 (n_19924, n_19918, n_19919);
  nand g47348 (n_20642, n_20634, n_20635);
  nand g47349 (n_19923, n_19916, n_19917);
  nand g47350 (n_20641, n_20632, n_20633);
  nand g47351 (n_19922, n_19914, n_19915);
  or g47352 (n_20712, wc452, n_16245);
  not gc452 (wc452, \data_stack_mem[4] [1]);
  or g47353 (n_22624, wc453, n_16127);
  not gc453 (wc453, \out_fifo[4][1] [8]);
  nand g47354 (n_19921, n_19912, n_19913);
  or g47355 (n_22627, wc454, n_16127);
  not gc454 (wc454, \out_fifo[4][1] [6]);
  or g47356 (n_18639, n_16110, n_16898);
  or g47357 (n_18640, wc455, n_16109);
  not gc455 (wc455, \out_fifo[7][2] [8]);
  or g47358 (n_18645, n_16113, n_16898);
  or g47359 (n_18646, wc456, n_16112);
  not gc456 (wc456, \out_fifo[5][2] [8]);
  or g47360 (n_18652, wc457, n_16115);
  not gc457 (wc457, \out_fifo[3][2] [8]);
  or g47361 (n_18657, n_16119, n_16898);
  or g47362 (n_18658, wc458, n_16118);
  not gc458 (wc458, \out_fifo[6][2] [8]);
  or g47363 (n_18663, n_16122, n_16898);
  or g47364 (n_18664, wc459, n_16121);
  not gc459 (wc459, \out_fifo[0][2] [8]);
  or g47365 (n_18669, n_16125, n_16898);
  or g47366 (n_18670, wc460, n_16124);
  not gc460 (wc460, \out_fifo[2][2] [8]);
  or g47367 (n_18675, n_16128, n_16898);
  or g47368 (n_18676, wc461, n_16127);
  not gc461 (wc461, \out_fifo[4][2] [8]);
  or g47369 (n_18681, n_16131, n_16898);
  or g47370 (n_18682, wc462, n_16130);
  not gc462 (wc462, \out_fifo[1][2] [8]);
  or g47371 (n_22630, wc463, n_16127);
  not gc463 (wc463, \out_fifo[4][1] [7]);
  or g47372 (n_18688, wc464, n_16109);
  not gc464 (wc464, \out_fifo[7][2] [0]);
  or g47373 (n_22633, wc465, n_16127);
  not gc465 (wc465, \out_fifo[4][1] [5]);
  or g47374 (n_22678, wc466, n_16109);
  not gc466 (wc466, \out_fifo[7][1] [1]);
  nand g47376 (n_19876, n_19870, n_19871);
  nand g47377 (n_19875, n_19868, n_19869);
  nand g47378 (n_18546, n_17303, n_16557);
  nand g47379 (n_19874, n_19866, n_19867);
  nand g47380 (n_19597, n_17429, n_19596);
  or g47381 (n_19040, n_19038, n_19039);
  or g47382 (n_22684, wc467, n_16112);
  not gc467 (wc467, \out_fifo[5][1] [1]);
  nand g47383 (n_24539, n_16506, n_16539);
  or g47384 (n_24540, n_16506, n_16539);
  nand g47385 (n_16540, n_24539, n_24540);
  nand g47386 (n_19873, n_19864, n_19865);
  nand g47387 (n_20596, n_20590, n_20591);
  or g47388 (n_22690, wc468, n_16115);
  not gc468 (wc468, \out_fifo[3][1] [1]);
  nand g47389 (n_20595, n_20588, n_20589);
  nand g47390 (n_20594, n_20586, n_20587);
  or g47391 (n_20700, wc469, n_16250);
  not gc469 (wc469, n_17640);
  nand g47392 (n_20593, n_20584, n_20585);
  or g47393 (n_20701, n_17640, wc470);
  not gc470 (wc470, n_16250);
  or g47394 (n_18694, wc471, n_16112);
  not gc471 (wc471, \out_fifo[5][2] [0]);
  or g47395 (n_22696, wc472, n_16118);
  not gc472 (wc472, \out_fifo[6][1] [1]);
  or g47396 (n_18700, wc473, n_16115);
  not gc473 (wc473, \out_fifo[3][2] [0]);
  or g47397 (n_22702, wc474, n_16121);
  not gc474 (wc474, \out_fifo[0][1] [1]);
  or g47398 (n_18706, wc475, n_16118);
  not gc475 (wc475, \out_fifo[6][2] [0]);
  or g47399 (n_22708, wc476, n_16124);
  not gc476 (wc476, \out_fifo[2][1] [1]);
  or g47400 (n_18712, wc477, n_16121);
  not gc477 (wc477, \out_fifo[0][2] [0]);
  or g47401 (n_22714, wc478, n_16127);
  not gc478 (wc478, \out_fifo[4][1] [1]);
  or g47402 (n_22720, wc479, n_16130);
  not gc479 (wc479, \out_fifo[1][1] [1]);
  or g47403 (n_18718, wc480, n_16124);
  not gc480 (wc480, \out_fifo[2][2] [0]);
  or g47404 (n_22726, wc481, n_16109);
  not gc481 (wc481, \out_fifo[7][1] [2]);
  or g47405 (n_18724, wc482, n_16127);
  not gc482 (wc482, \out_fifo[4][2] [0]);
  or g47406 (n_22732, wc483, n_16112);
  not gc483 (wc483, \out_fifo[5][1] [2]);
  or g47407 (n_18730, wc484, n_16130);
  not gc484 (wc484, \out_fifo[1][2] [0]);
  or g47408 (n_22738, wc485, n_16115);
  not gc485 (wc485, \out_fifo[3][1] [2]);
  or g47409 (n_18735, n_16110, n_16143);
  or g47410 (n_18736, wc486, n_16109);
  not gc486 (wc486, \out_fifo[7][2] [1]);
  or g47411 (n_22744, wc487, n_16118);
  not gc487 (wc487, \out_fifo[6][1] [2]);
  or g47412 (n_18741, n_16113, n_16143);
  or g47413 (n_18742, wc488, n_16112);
  not gc488 (wc488, \out_fifo[5][2] [1]);
  or g47414 (n_18748, wc489, n_16115);
  not gc489 (wc489, \out_fifo[3][2] [1]);
  or g47415 (n_18753, n_16119, n_16143);
  or g47416 (n_18754, wc490, n_16118);
  not gc490 (wc490, \out_fifo[6][2] [1]);
  or g47417 (n_18759, n_16122, n_16143);
  or g47418 (n_18760, wc491, n_16121);
  not gc491 (wc491, \out_fifo[0][2] [1]);
  or g47419 (n_18765, n_16125, n_16143);
  or g47420 (n_18766, wc492, n_16124);
  not gc492 (wc492, \out_fifo[2][2] [1]);
  or g47421 (n_18771, n_16128, n_16143);
  or g47422 (n_18772, wc493, n_16127);
  not gc493 (wc493, \out_fifo[4][2] [1]);
  or g47423 (n_18777, n_16131, n_16143);
  or g47424 (n_18778, wc494, n_16130);
  not gc494 (wc494, \out_fifo[1][2] [1]);
  nand g47425 (n_19828, n_19822, n_19823);
  nand g47426 (n_19827, n_19820, n_19821);
  nand g47427 (n_19826, n_19818, n_19819);
  nand g47428 (n_19825, n_19816, n_19817);
  or g47429 (n_22750, wc495, n_16121);
  not gc495 (wc495, \out_fifo[0][1] [2]);
  nand g47430 (n_19780, n_19774, n_19775);
  nand g47431 (n_19779, n_19772, n_19773);
  nand g47432 (n_19778, n_19770, n_19771);
  nand g47433 (n_20161, n_20152, n_20153);
  nand g47434 (n_19777, n_19768, n_19769);
  or g47435 (n_22756, wc496, n_16124);
  not gc496 (wc496, \out_fifo[2][1] [2]);
  nand g47436 (n_20548, n_20542, n_20543);
  nand g47437 (n_20547, n_20540, n_20541);
  nand g47438 (n_20546, n_20538, n_20539);
  nand g47439 (n_20545, n_20536, n_20537);
  nand g47440 (n_19732, n_19726, n_19727);
  nand g47441 (n_19731, n_19724, n_19725);
  nand g47442 (n_18325, n_18323, n_18324);
  nand g47443 (n_19730, n_19722, n_19723);
  nand g47444 (n_19729, n_19720, n_19721);
  nand g47445 (n_22993, n_17425, n_16523);
  or g47446 (n_22762, wc497, n_16127);
  not gc497 (wc497, \out_fifo[4][1] [2]);
  or g47447 (n_20706, \data_stack_mem[4] [1], wc498);
  not gc498 (wc498, n_16220);
  nand g47448 (n_19684, n_19678, n_19679);
  nand g47449 (n_19683, n_19676, n_19677);
  nand g47450 (n_20162, n_20154, n_20155);
  nand g47451 (n_19682, n_19674, n_19675);
  nand g47452 (n_19681, n_19672, n_19673);
  nand g47453 (n_20500, n_20494, n_20495);
  nand g47454 (n_20499, n_20492, n_20493);
  nand g47455 (n_20353, n_20344, n_20345);
  nand g47456 (n_20498, n_20490, n_20491);
  nand g47457 (n_20497, n_20488, n_20489);
  nand g47458 (n_19637, n_19632, n_19633);
  nand g47459 (n_19636, n_19630, n_19631);
  nand g47460 (n_19635, n_19628, n_19629);
  nand g47461 (n_19634, n_19626, n_19627);
  or g47462 (n_22768, wc499, n_16130);
  not gc499 (wc499, \out_fifo[1][1] [2]);
  or g47463 (n_22780, wc500, n_16109);
  not gc500 (wc500, \out_fifo[7][0] [0]);
  or g47464 (n_22786, wc501, n_16112);
  not gc501 (wc501, \out_fifo[5][0] [0]);
  nand g47465 (n_20163, n_20156, n_20157);
  or g47466 (n_19100, n_19098, n_19099);
  nand g47467 (n_20452, n_20446, n_20447);
  nand g47468 (n_20451, n_20444, n_20445);
  nand g47469 (n_20450, n_20442, n_20443);
  or g47470 (n_17009, wc502, n_16986);
  not gc502 (wc502, n_19105);
  nand g47471 (n_20449, n_20440, n_20441);
  or g47473 (n_22792, wc503, n_16115);
  not gc503 (wc503, \out_fifo[3][0] [0]);
  nand g47476 (n_16282, n_24541, n_24542);
  nand g47477 (n_24543, n_16366, n_16367);
  or g47478 (n_24544, n_16366, n_16367);
  nand g47479 (n_16368, n_24543, n_24544);
  nand g47481 (n_20164, n_20158, n_20159);
  nand g47484 (n_20354, n_20346, n_20347);
  or g47485 (n_22798, wc504, n_16118);
  not gc504 (wc504, \out_fifo[6][0] [0]);
  or g47486 (n_22804, wc505, n_16121);
  not gc505 (wc505, \out_fifo[0][0] [0]);
  or g47487 (n_22810, wc506, n_16124);
  not gc506 (wc506, \out_fifo[2][0] [0]);
  or g47488 (n_22816, wc507, n_16127);
  not gc507 (wc507, \out_fifo[4][0] [0]);
  or g47489 (n_18538, n_16522, n_16523);
  or g47490 (n_22822, wc508, n_16130);
  not gc508 (wc508, \out_fifo[1][0] [0]);
  or g47491 (n_22843, wc509, n_16109);
  not gc509 (wc509, \out_fifo[7][1] [3]);
  or g47492 (n_22849, wc510, n_16112);
  not gc510 (wc510, \out_fifo[5][1] [3]);
  or g47493 (n_22855, wc511, n_16115);
  not gc511 (wc511, \out_fifo[3][1] [3]);
  nand g47494 (n_20355, n_20348, n_20349);
  or g47495 (n_22861, wc512, n_16118);
  not gc512 (wc512, \out_fifo[6][1] [3]);
  nand g47496 (n_20356, n_20350, n_20351);
  or g47497 (n_22867, wc513, n_16121);
  not gc513 (wc513, \out_fifo[0][1] [3]);
  or g47498 (n_22873, wc514, n_16124);
  not gc514 (wc514, \out_fifo[2][1] [3]);
  nand g47501 (n_16211, n_24545, n_24546);
  nand g47502 (n_18537, n_16521, n_16523);
  or g47503 (n_22879, wc515, n_16127);
  not gc515 (wc515, \out_fifo[4][1] [3]);
  or g47504 (n_22885, wc516, n_16130);
  not gc516 (wc516, \out_fifo[1][1] [3]);
  or g47505 (n_22891, wc517, n_16109);
  not gc517 (wc517, \out_fifo[7][1] [4]);
  or g47506 (n_22897, wc518, n_16112);
  not gc518 (wc518, \out_fifo[5][1] [4]);
  or g47507 (n_22903, wc519, n_16115);
  not gc519 (wc519, \out_fifo[3][1] [4]);
  or g47508 (n_22909, wc520, n_16118);
  not gc520 (wc520, \out_fifo[6][1] [4]);
  nand g47509 (n_20404, n_20398, n_20399);
  nand g47510 (n_20403, n_20396, n_20397);
  nand g47511 (n_24547, n_16155, n_16167);
  or g47512 (n_24548, n_16155, n_16167);
  nand g47513 (n_16168, n_24547, n_24548);
  nand g47514 (n_20402, n_20394, n_20395);
  nand g47515 (n_20209, n_20200, n_20201);
  nand g47516 (n_20401, n_20392, n_20393);
  or g47517 (n_22915, wc521, n_16121);
  not gc521 (wc521, \out_fifo[0][1] [4]);
  nand g47518 (n_20210, n_20202, n_20203);
  nand g47519 (n_20211, n_20204, n_20205);
  nand g47520 (n_20212, n_20206, n_20207);
  nand g47521 (n_24549, n_17390, n_16108);
  or g47522 (n_24550, n_17390, n_16108);
  nand g47523 (n_16907, n_24549, n_24550);
  or g47524 (n_22921, wc522, n_16124);
  not gc522 (wc522, \out_fifo[2][1] [4]);
  or g47525 (n_22927, wc523, n_16127);
  not gc523 (wc523, \out_fifo[4][1] [4]);
  or g47526 (n_22933, wc524, n_16130);
  not gc524 (wc524, \out_fifo[1][1] [4]);
  nand g47527 (n_18349, n_18347, n_18348);
  or g47528 (n_22939, wc525, n_16109);
  not gc525 (wc525, \out_fifo[7][1] [0]);
  or g47529 (n_22945, wc526, n_16112);
  not gc526 (wc526, \out_fifo[5][1] [0]);
  or g47530 (n_22951, wc527, n_16115);
  not gc527 (wc527, \out_fifo[3][1] [0]);
  nand g47531 (n_20257, n_20248, n_20249);
  or g47532 (n_22957, wc528, n_16118);
  not gc528 (wc528, \out_fifo[6][1] [0]);
  or g47533 (n_22963, wc529, n_16121);
  not gc529 (wc529, \out_fifo[0][1] [0]);
  or g47534 (n_22969, wc530, n_16124);
  not gc530 (wc530, \out_fifo[2][1] [0]);
  or g47535 (n_22975, wc531, n_16127);
  not gc531 (wc531, \out_fifo[4][1] [0]);
  or g47536 (n_22981, wc532, n_16130);
  not gc532 (wc532, \out_fifo[1][1] [0]);
  nand g47537 (n_20258, n_20250, n_20251);
  nand g47538 (n_17061, n_23022, n_23023);
  nand g47540 (n_20259, n_20252, n_20253);
  nand g47541 (n_20260, n_20254, n_20255);
  or g47543 (n_20394, wc533, n_17077);
  not gc533 (wc533, \out_fifo[1][0] [6]);
  or g47545 (n_19359, wc534, n_16997);
  not gc534 (wc534, sh_reg_in[2]);
  or g47546 (n_19353, wc535, n_16997);
  not gc535 (wc535, sh_reg_in[6]);
  or g47547 (n_19347, wc536, n_16997);
  not gc536 (wc536, sh_reg_in[0]);
  or g47548 (n_20393, wc537, n_17079);
  not gc537 (wc537, \out_fifo[5][0] [6]);
  or g47549 (n_19341, wc538, n_16997);
  not gc538 (wc538, sh_reg_in[4]);
  or g47550 (n_19335, wc539, n_16997);
  not gc539 (wc539, sh_reg_in[7]);
  or g47551 (n_19329, wc540, n_16997);
  not gc540 (wc540, sh_reg_in[5]);
  or g47552 (n_19323, wc541, n_16997);
  not gc541 (wc541, sh_reg_in[1]);
  or g47553 (n_19317, wc542, n_16997);
  not gc542 (wc542, sh_reg_in[3]);
  or g47554 (n_20392, wc543, n_17078);
  not gc543 (wc543, \out_fifo[4][0] [6]);
  or g47556 (n_20395, wc544, n_17076);
  not gc544 (wc544, \out_fifo[0][0] [6]);
  or g47557 (n_20397, wc545, n_17068);
  not gc545 (wc545, \out_fifo[7][0] [6]);
  or g47558 (n_20398, wc546, n_17070);
  not gc546 (wc546, \out_fifo[2][0] [6]);
  or g47559 (n_20399, wc547, n_17072);
  not gc547 (wc547, \out_fifo[3][0] [6]);
  or g47560 (n_20400, wc548, n_17074);
  not gc548 (wc548, \out_fifo[6][0] [6]);
  or g47562 (n_19251, wc549, n_16962);
  not gc549 (wc549, sh_reg_in[2]);
  or g47563 (n_19245, wc550, n_16962);
  not gc550 (wc550, sh_reg_in[0]);
  or g47564 (n_19239, wc551, n_16962);
  not gc551 (wc551, sh_reg_in[4]);
  or g47565 (n_19233, wc552, n_16962);
  not gc552 (wc552, sh_reg_in[5]);
  or g47566 (n_19227, wc553, n_16962);
  not gc553 (wc553, sh_reg_in[6]);
  or g47567 (n_19221, wc554, n_16962);
  not gc554 (wc554, sh_reg_in[7]);
  or g47568 (n_19215, wc555, n_16962);
  not gc555 (wc555, sh_reg_in[1]);
  or g47569 (n_19209, wc556, n_16962);
  not gc556 (wc556, sh_reg_in[3]);
  or g47571 (n_19197, wc557, n_16950);
  not gc557 (wc557, sh_reg_in[7]);
  or g47572 (n_19191, wc558, n_16950);
  not gc558 (wc558, sh_reg_in[0]);
  or g47573 (n_19482, wc559, n_17008);
  not gc559 (wc559, sh_reg_in[2]);
  or g47574 (n_19185, wc560, n_16950);
  not gc560 (wc560, sh_reg_in[6]);
  or g47575 (n_19488, wc561, n_17008);
  not gc561 (wc561, sh_reg_in[0]);
  or g47576 (n_19179, wc562, n_16950);
  not gc562 (wc562, sh_reg_in[4]);
  or g47577 (n_19494, wc563, n_17008);
  not gc563 (wc563, sh_reg_in[7]);
  or g47578 (n_19173, wc564, n_16950);
  not gc564 (wc564, sh_reg_in[3]);
  or g47579 (n_19500, wc565, n_17008);
  not gc565 (wc565, sh_reg_in[5]);
  or g47580 (n_19167, wc566, n_16950);
  not gc566 (wc566, sh_reg_in[1]);
  or g47581 (n_19506, wc567, n_17008);
  not gc567 (wc567, n_16946);
  or g47582 (n_20440, wc568, n_17078);
  not gc568 (wc568, \out_fifo[4][0] [7]);
  or g47583 (n_19512, wc569, n_17008);
  not gc569 (wc569, sh_reg_in[4]);
  or g47584 (n_20441, wc570, n_17079);
  not gc570 (wc570, \out_fifo[5][0] [7]);
  or g47585 (n_19518, wc571, n_17008);
  not gc571 (wc571, sh_reg_in[3]);
  or g47586 (n_20442, wc572, n_17077);
  not gc572 (wc572, \out_fifo[1][0] [7]);
  nand g47589 (n_16784, n_24551, n_24552);
  or g47590 (n_19524, wc573, n_17008);
  not gc573 (wc573, sh_reg_in[1]);
  or g47591 (n_19161, wc574, n_16950);
  not gc574 (wc574, sh_reg_in[2]);
  or g47592 (n_19530, wc575, n_17008);
  not gc575 (wc575, sh_reg_in[6]);
  or g47593 (n_19155, wc576, n_16950);
  not gc576 (wc576, sh_reg_in[5]);
  or g47594 (n_19536, wc577, n_17020);
  not gc577 (wc577, sh_reg_in[0]);
  or g47595 (n_20443, wc578, n_17076);
  not gc578 (wc578, \out_fifo[0][0] [7]);
  nand g47598 (n_16280, n_24553, n_24554);
  or g47599 (n_19542, wc579, n_17020);
  not gc579 (wc579, sh_reg_in[1]);
  or g47600 (n_20445, wc580, n_17068);
  not gc580 (wc580, \out_fifo[7][0] [7]);
  nand g47601 (n_19144, n_19142, n_19143);
  or g47602 (n_19548, wc581, n_17020);
  not gc581 (wc581, sh_reg_in[2]);
  or g47603 (n_20446, wc582, n_17070);
  not gc582 (wc582, \out_fifo[2][0] [7]);
  or g47604 (n_20447, wc583, n_17072);
  not gc583 (wc583, \out_fifo[3][0] [7]);
  or g47605 (n_19554, wc584, n_17020);
  not gc584 (wc584, sh_reg_in[3]);
  or g47606 (n_20448, wc585, n_17074);
  not gc585 (wc585, \out_fifo[6][0] [7]);
  or g47607 (n_19560, wc586, n_17020);
  not gc586 (wc586, sh_reg_in[5]);
  or g47609 (n_19566, wc587, n_17020);
  not gc587 (wc587, sh_reg_in[6]);
  or g47610 (n_20488, wc588, n_17078);
  not gc588 (wc588, \out_fifo[4][0] [8]);
  or g47611 (n_19572, wc589, n_17020);
  not gc589 (wc589, sh_reg_in[7]);
  or g47612 (n_20489, wc590, n_17079);
  not gc590 (wc590, \out_fifo[5][0] [8]);
  or g47613 (n_19578, wc591, n_17020);
  not gc591 (wc591, n_16946);
  nand g47614 (n_16983, n_18891, n_18892);
  or g47615 (n_19584, wc592, n_17020);
  not gc592 (wc592, sh_reg_in[4]);
  or g47616 (n_20490, wc593, n_17077);
  not gc593 (wc593, \out_fifo[1][0] [8]);
  or g47617 (n_19626, wc594, n_17079);
  not gc594 (wc594, \out_fifo[5][0] [0]);
  or g47618 (n_19627, wc595, n_17078);
  not gc595 (wc595, \out_fifo[4][0] [0]);
  or g47619 (n_19628, wc596, n_17077);
  not gc596 (wc596, \out_fifo[1][0] [0]);
  or g47620 (n_19629, wc597, n_17076);
  not gc597 (wc597, \out_fifo[0][0] [0]);
  or g47621 (n_19630, wc598, n_17074);
  not gc598 (wc598, \out_fifo[6][0] [0]);
  or g47622 (n_19631, wc599, n_17072);
  not gc599 (wc599, \out_fifo[3][0] [0]);
  or g47623 (n_19632, wc600, n_17070);
  not gc600 (wc600, \out_fifo[2][0] [0]);
  or g47624 (n_19633, wc601, n_17068);
  not gc601 (wc601, \out_fifo[7][0] [0]);
  or g47625 (n_20491, wc602, n_17076);
  not gc602 (wc602, \out_fifo[0][0] [8]);
  nand g47626 (n_16982, n_18885, n_18886);
  or g47627 (n_20493, wc603, n_17068);
  not gc603 (wc603, \out_fifo[7][0] [8]);
  or g47628 (n_20494, wc604, n_17070);
  not gc604 (wc604, \out_fifo[2][0] [8]);
  nand g47629 (n_16981, n_18879, n_18880);
  or g47630 (n_20495, wc605, n_17072);
  not gc605 (wc605, \out_fifo[3][0] [8]);
  or g47631 (n_20496, wc606, n_17074);
  not gc606 (wc606, \out_fifo[6][0] [8]);
  or g47632 (n_19672, wc607, n_17078);
  not gc607 (wc607, \out_fifo[4][1] [1]);
  or g47633 (n_19673, wc608, n_17079);
  not gc608 (wc608, \out_fifo[5][1] [1]);
  or g47634 (n_19674, wc609, n_17077);
  not gc609 (wc609, \out_fifo[1][1] [1]);
  or g47635 (n_19675, wc610, n_17076);
  not gc610 (wc610, \out_fifo[0][1] [1]);
  nand g47636 (n_16980, n_18873, n_18874);
  or g47637 (n_19677, wc611, n_17068);
  not gc611 (wc611, \out_fifo[7][1] [1]);
  or g47638 (n_19678, wc612, n_17070);
  not gc612 (wc612, \out_fifo[2][1] [1]);
  or g47639 (n_19679, wc613, n_17072);
  not gc613 (wc613, \out_fifo[3][1] [1]);
  or g47640 (n_19680, wc614, n_17074);
  not gc614 (wc614, \out_fifo[6][1] [1]);
  nand g47641 (n_16979, n_18867, n_18868);
  nand g47642 (n_16978, n_18861, n_18862);
  nand g47643 (n_16977, n_18855, n_18856);
  or g47644 (n_20536, wc615, n_17078);
  not gc615 (wc615, \out_fifo[4][2] [1]);
  nand g47645 (n_16976, n_18849, n_18850);
  or g47646 (n_20537, wc616, n_17079);
  not gc616 (wc616, \out_fifo[5][2] [1]);
  or g47647 (n_20538, wc617, n_17077);
  not gc617 (wc617, \out_fifo[1][2] [1]);
  nand g47648 (n_16975, n_18843, n_18844);
  or g47649 (n_20539, wc618, n_17076);
  not gc618 (wc618, \out_fifo[0][2] [1]);
  or g47650 (n_20541, wc619, n_17068);
  not gc619 (wc619, \out_fifo[7][2] [1]);
  nand g47651 (n_17052, n_18837, n_18838);
  or g47652 (n_19720, wc620, n_17078);
  not gc620 (wc620, \out_fifo[4][1] [3]);
  or g47653 (n_19721, wc621, n_17079);
  not gc621 (wc621, \out_fifo[5][1] [3]);
  or g47654 (n_19722, wc622, n_17077);
  not gc622 (wc622, \out_fifo[1][1] [3]);
  or g47655 (n_19723, wc623, n_17076);
  not gc623 (wc623, \out_fifo[0][1] [3]);
  or g47656 (n_20352, wc624, n_17074);
  not gc624 (wc624, \out_fifo[6][0] [5]);
  or g47657 (n_19725, wc625, n_17068);
  not gc625 (wc625, \out_fifo[7][1] [3]);
  or g47658 (n_19726, wc626, n_17070);
  not gc626 (wc626, \out_fifo[2][1] [3]);
  or g47659 (n_19727, wc627, n_17072);
  not gc627 (wc627, \out_fifo[3][1] [3]);
  or g47660 (n_19728, wc628, n_17074);
  not gc628 (wc628, \out_fifo[6][1] [3]);
  or g47661 (n_20542, wc629, n_17070);
  not gc629 (wc629, \out_fifo[2][2] [1]);
  or g47662 (n_20543, wc630, n_17072);
  not gc630 (wc630, \out_fifo[3][2] [1]);
  nand g47663 (n_16947, n_18831, n_18832);
  nand g47664 (n_16938, n_18825, n_18826);
  or g47666 (n_20544, wc631, n_17074);
  not gc631 (wc631, \out_fifo[6][2] [1]);
  nand g47667 (n_16937, n_18819, n_18820);
  or g47668 (n_19768, wc632, n_17078);
  not gc632 (wc632, \out_fifo[4][1] [4]);
  or g47669 (n_19769, wc633, n_17079);
  not gc633 (wc633, \out_fifo[5][1] [4]);
  or g47670 (n_19770, wc634, n_17077);
  not gc634 (wc634, \out_fifo[1][1] [4]);
  or g47671 (n_19771, wc635, n_17076);
  not gc635 (wc635, \out_fifo[0][1] [4]);
  or g47672 (n_20351, wc636, n_17072);
  not gc636 (wc636, \out_fifo[3][0] [5]);
  or g47673 (n_19773, wc637, n_17068);
  not gc637 (wc637, \out_fifo[7][1] [4]);
  or g47674 (n_19774, wc638, n_17070);
  not gc638 (wc638, \out_fifo[2][1] [4]);
  or g47675 (n_19775, wc639, n_17072);
  not gc639 (wc639, \out_fifo[3][1] [4]);
  or g47676 (n_19776, wc640, n_17074);
  not gc640 (wc640, \out_fifo[6][1] [4]);
  nand g47677 (n_16935, n_18807, n_18808);
  nand g47678 (n_16934, n_18801, n_18802);
  or g47679 (n_20584, wc641, n_17072);
  not gc641 (wc641, \out_fifo[3][2] [6]);
  nand g47680 (n_16933, n_18795, n_18796);
  or g47681 (n_20585, wc642, n_17070);
  not gc642 (wc642, \out_fifo[2][2] [6]);
  or g47682 (n_20586, wc643, n_17068);
  not gc643 (wc643, \out_fifo[7][2] [6]);
  nand g47683 (n_16932, n_18789, n_18790);
  or g47684 (n_19816, wc644, n_17078);
  not gc644 (wc644, \out_fifo[4][1] [5]);
  or g47685 (n_19817, wc645, n_17079);
  not gc645 (wc645, \out_fifo[5][1] [5]);
  or g47686 (n_19818, wc646, n_17077);
  not gc646 (wc646, \out_fifo[1][1] [5]);
  or g47687 (n_19819, wc647, n_17076);
  not gc647 (wc647, \out_fifo[0][1] [5]);
  or g47688 (n_20350, wc648, n_17070);
  not gc648 (wc648, \out_fifo[2][0] [5]);
  or g47689 (n_19821, wc649, n_17068);
  not gc649 (wc649, \out_fifo[7][1] [5]);
  or g47690 (n_19822, wc650, n_17070);
  not gc650 (wc650, \out_fifo[2][1] [5]);
  or g47691 (n_19823, wc651, n_17072);
  not gc651 (wc651, \out_fifo[3][1] [5]);
  or g47692 (n_19824, wc652, n_17074);
  not gc652 (wc652, \out_fifo[6][1] [5]);
  or g47693 (n_20587, wc653, n_17074);
  not gc653 (wc653, \out_fifo[6][2] [6]);
  or g47694 (n_20589, wc654, n_17076);
  not gc654 (wc654, \out_fifo[0][2] [6]);
  nand g47695 (n_16931, n_18783, n_18784);
  or g47696 (n_20590, wc655, n_17077);
  not gc655 (wc655, \out_fifo[1][2] [6]);
  or g47697 (n_20591, wc656, n_17078);
  not gc656 (wc656, \out_fifo[4][2] [6]);
  or g47698 (n_18747, n_16116, n_16143);
  or g47699 (n_20592, wc657, n_17079);
  not gc657 (wc657, \out_fifo[5][2] [6]);
  or g47700 (n_19864, wc658, n_17078);
  not gc658 (wc658, \out_fifo[4][1] [2]);
  or g47701 (n_19865, wc659, n_17079);
  not gc659 (wc659, \out_fifo[5][1] [2]);
  or g47702 (n_19866, wc660, n_17077);
  not gc660 (wc660, \out_fifo[1][1] [2]);
  or g47703 (n_19867, wc661, n_17076);
  not gc661 (wc661, \out_fifo[0][1] [2]);
  or g47704 (n_20349, wc662, n_17068);
  not gc662 (wc662, \out_fifo[7][0] [5]);
  or g47705 (n_19869, wc663, n_17068);
  not gc663 (wc663, \out_fifo[7][1] [2]);
  or g47706 (n_19870, wc664, n_17070);
  not gc664 (wc664, \out_fifo[2][1] [2]);
  or g47707 (n_19871, wc665, n_17072);
  not gc665 (wc665, \out_fifo[3][1] [2]);
  or g47708 (n_19872, wc666, n_17074);
  not gc666 (wc666, \out_fifo[6][1] [2]);
  nand g47709 (n_17640, n_18903, n_18904);
  or g47710 (n_20632, wc667, n_17072);
  not gc667 (wc667, \out_fifo[3][0] [2]);
  or g47711 (n_20633, wc668, n_17070);
  not gc668 (wc668, \out_fifo[2][0] [2]);
  or g47712 (n_19039, wc669, n_19037);
  not gc669 (wc669, n_19036);
  or g47713 (n_20634, wc670, n_17068);
  not gc670 (wc670, \out_fifo[7][0] [2]);
  or g47714 (n_19596, wc671, n_16247);
  not gc671 (wc671, \data_stack_mem[3] [1]);
  or g47715 (n_20635, wc672, n_17074);
  not gc672 (wc672, \out_fifo[6][0] [2]);
  or g47716 (n_20637, wc673, n_17076);
  not gc673 (wc673, \out_fifo[0][0] [2]);
  or g47717 (n_20638, wc674, n_17077);
  not gc674 (wc674, \out_fifo[1][0] [2]);
  or g47719 (n_18651, n_16116, n_16898);
  or g47720 (n_19912, wc675, n_17078);
  not gc675 (wc675, \out_fifo[4][1] [7]);
  or g47721 (n_19913, wc676, n_17079);
  not gc676 (wc676, \out_fifo[5][1] [7]);
  or g47722 (n_19914, wc677, n_17077);
  not gc677 (wc677, \out_fifo[1][1] [7]);
  or g47723 (n_19915, wc678, n_17076);
  not gc678 (wc678, \out_fifo[0][1] [7]);
  or g47724 (n_20347, wc679, n_17076);
  not gc679 (wc679, \out_fifo[0][0] [5]);
  or g47725 (n_19917, wc680, n_17068);
  not gc680 (wc680, \out_fifo[7][1] [7]);
  or g47726 (n_19918, wc681, n_17070);
  not gc681 (wc681, \out_fifo[2][1] [7]);
  or g47727 (n_19919, wc682, n_17072);
  not gc682 (wc682, \out_fifo[3][1] [7]);
  or g47728 (n_19920, wc683, n_17074);
  not gc683 (wc683, \out_fifo[6][1] [7]);
  or g47729 (n_20639, wc684, n_17078);
  not gc684 (wc684, \out_fifo[4][0] [2]);
  or g47730 (n_20640, wc685, n_17079);
  not gc685 (wc685, \out_fifo[5][0] [2]);
  or g47731 (n_19009, wc686, n_19007);
  not gc686 (wc686, n_19006);
  or g47733 (n_20680, wc687, n_17072);
  not gc687 (wc687, \out_fifo[3][0] [3]);
  or g47734 (n_19960, wc688, n_17078);
  not gc688 (wc688, \out_fifo[4][1] [8]);
  or g47735 (n_19961, wc689, n_17079);
  not gc689 (wc689, \out_fifo[5][1] [8]);
  or g47736 (n_19962, wc690, n_17077);
  not gc690 (wc690, \out_fifo[1][1] [8]);
  or g47737 (n_19963, wc691, n_17076);
  not gc691 (wc691, \out_fifo[0][1] [8]);
  or g47738 (n_20346, wc692, n_17077);
  not gc692 (wc692, \out_fifo[1][0] [5]);
  or g47739 (n_19965, wc693, n_17068);
  not gc693 (wc693, \out_fifo[7][1] [8]);
  or g47740 (n_19966, wc694, n_17070);
  not gc694 (wc694, \out_fifo[2][1] [8]);
  or g47741 (n_19967, wc695, n_17072);
  not gc695 (wc695, \out_fifo[3][1] [8]);
  or g47742 (n_19968, wc696, n_17074);
  not gc696 (wc696, \out_fifo[6][1] [8]);
  or g47743 (n_20681, wc697, n_17070);
  not gc697 (wc697, \out_fifo[2][0] [3]);
  or g47744 (n_20682, wc698, n_17068);
  not gc698 (wc698, \out_fifo[7][0] [3]);
  or g47746 (n_20683, wc699, n_17074);
  not gc699 (wc699, \out_fifo[6][0] [3]);
  nand g47749 (n_16445, n_24555, n_24556);
  or g47750 (n_20685, wc700, n_17076);
  not gc700 (wc700, \out_fifo[0][0] [3]);
  or g47751 (n_20686, wc701, n_17077);
  not gc701 (wc701, \out_fifo[1][0] [3]);
  nand g47754 (n_16602, n_24557, n_24558);
  or g47756 (n_20345, wc702, n_17079);
  not gc702 (wc702, \out_fifo[5][0] [5]);
  or g47757 (n_20344, wc703, n_17078);
  not gc703 (wc703, \out_fifo[4][0] [5]);
  or g47758 (n_20687, wc704, n_17078);
  not gc704 (wc704, \out_fifo[4][0] [3]);
  or g47759 (n_20008, wc705, n_17078);
  not gc705 (wc705, \out_fifo[4][2] [8]);
  or g47760 (n_20009, wc706, n_17079);
  not gc706 (wc706, \out_fifo[5][2] [8]);
  or g47761 (n_20010, wc707, n_17077);
  not gc707 (wc707, \out_fifo[1][2] [8]);
  or g47762 (n_20011, wc708, n_17076);
  not gc708 (wc708, \out_fifo[0][2] [8]);
  or g47763 (n_20688, wc709, n_17079);
  not gc709 (wc709, \out_fifo[5][0] [3]);
  or g47764 (n_20013, wc710, n_17068);
  not gc710 (wc710, \out_fifo[7][2] [8]);
  nand g47765 (n_18559, n_18557, n_18558);
  or g47766 (n_20014, wc711, n_17070);
  not gc711 (wc711, \out_fifo[2][2] [8]);
  or g47767 (n_20015, wc712, n_17072);
  not gc712 (wc712, \out_fifo[3][2] [8]);
  or g47768 (n_20016, wc713, n_17074);
  not gc713 (wc713, \out_fifo[6][2] [8]);
  or g47769 (n_19069, wc714, n_19067);
  not gc714 (wc714, n_19066);
  or g47771 (n_19471, \data_stack_mem[2] [1], wc715);
  not gc715 (wc715, n_16226);
  nand g47772 (n_17058, n_18465, n_18466);
  nand g47773 (n_16925, n_18456, n_18457);
  nand g47774 (n_17060, n_18444, n_18445);
  nand g47776 (n_17051, n_18435, n_18436);
  nand g47777 (n_17050, n_18429, n_18430);
  nand g47778 (n_17049, n_18423, n_18424);
  or g47779 (n_18980, n_18977, n_18978);
  nand g47780 (n_17048, n_18417, n_18418);
  nand g47782 (n_16557, n_18151, n_23008);
  nand g47783 (n_17047, n_18411, n_18412);
  nand g47784 (n_17046, n_18405, n_18406);
  nand g47785 (n_17045, n_18399, n_18400);
  or g47786 (n_20056, wc716, n_17078);
  not gc716 (wc716, \out_fifo[4][2] [9]);
  or g47787 (n_20057, wc717, n_17079);
  not gc717 (wc717, \out_fifo[5][2] [9]);
  or g47788 (n_20058, wc718, n_17077);
  not gc718 (wc718, \out_fifo[1][2] [9]);
  or g47789 (n_20059, wc719, n_17076);
  not gc719 (wc719, \out_fifo[0][2] [9]);
  nand g47790 (n_17044, n_18393, n_18394);
  or g47791 (n_20061, wc720, n_17068);
  not gc720 (wc720, \out_fifo[7][2] [9]);
  or g47792 (n_20062, wc721, n_17070);
  not gc721 (wc721, \out_fifo[2][2] [9]);
  or g47793 (n_20063, wc722, n_17072);
  not gc722 (wc722, \out_fifo[3][2] [9]);
  or g47794 (n_20064, wc723, n_17074);
  not gc723 (wc723, \out_fifo[6][2] [9]);
  or g47795 (n_19463, n_16224, n_16226);
  or g47796 (n_18946, wc724, n_18944);
  not gc724 (wc724, n_18943);
  nand g47799 (n_18913, n_18911, n_18912);
  or g47800 (n_19590, \data_stack_mem[3] [1], wc725);
  not gc725 (wc725, n_16222);
  or g47801 (n_20104, wc726, n_17078);
  not gc726 (wc726, \out_fifo[4][1] [6]);
  or g47802 (n_20105, wc727, n_17079);
  not gc727 (wc727, \out_fifo[5][1] [6]);
  or g47803 (n_20106, wc728, n_17077);
  not gc728 (wc728, \out_fifo[1][1] [6]);
  or g47804 (n_20107, wc729, n_17076);
  not gc729 (wc729, \out_fifo[0][1] [6]);
  or g47805 (n_18034, n_18033, n_16179);
  or g47806 (n_20109, wc730, n_17068);
  not gc730 (wc730, \out_fifo[7][1] [6]);
  or g47807 (n_20110, wc731, n_17070);
  not gc731 (wc731, \out_fifo[2][1] [6]);
  or g47808 (n_20111, wc732, n_17072);
  not gc732 (wc732, \out_fifo[3][1] [6]);
  or g47809 (n_20112, wc733, n_17074);
  not gc733 (wc733, \out_fifo[6][1] [6]);
  or g47811 (n_18103, n_18101, wc734);
  not gc734 (wc734, rst_n);
  nand g47813 (n_17056, n_17964, n_17965);
  or g47814 (n_20152, wc735, n_17078);
  not gc735 (wc735, \out_fifo[4][2] [0]);
  or g47815 (n_20153, wc736, n_17079);
  not gc736 (wc736, \out_fifo[5][2] [0]);
  or g47816 (n_20154, wc737, n_17077);
  not gc737 (wc737, \out_fifo[1][2] [0]);
  or g47817 (n_20155, wc738, n_17076);
  not gc738 (wc738, \out_fifo[0][2] [0]);
  or g47818 (n_20304, wc739, n_17074);
  not gc739 (wc739, \out_fifo[6][0] [4]);
  or g47819 (n_20157, wc740, n_17068);
  not gc740 (wc740, \out_fifo[7][2] [0]);
  or g47820 (n_20158, wc741, n_17070);
  not gc741 (wc741, \out_fifo[2][2] [0]);
  or g47821 (n_20159, wc742, n_17072);
  not gc742 (wc742, \out_fifo[3][2] [0]);
  or g47822 (n_20160, wc743, n_17074);
  not gc743 (wc743, \out_fifo[6][2] [0]);
  nand g47823 (n_24559, n_16502, n_16538);
  or g47824 (n_24560, n_16502, n_16538);
  nand g47825 (n_16539, n_24559, n_24560);
  or g47826 (n_20303, wc744, n_17072);
  not gc744 (wc744, \out_fifo[3][0] [4]);
  or g47827 (n_20302, wc745, n_17070);
  not gc745 (wc745, \out_fifo[2][0] [4]);
  or g47828 (n_20301, wc746, n_17068);
  not gc746 (wc746, \out_fifo[7][0] [4]);
  or g47831 (n_19099, wc747, n_19097);
  not gc747 (wc747, n_19096);
  nand g47833 (n_24562, n_16355, n_16365);
  or g47834 (n_24563, n_16355, n_16365);
  nand g47835 (n_16366, n_24562, n_24563);
  nand g47836 (n_16109, rst_n, n_16079);
  or g47837 (n_16110, n_16079, wc748);
  not gc748 (wc748, rst_n);
  nand g47838 (n_16112, rst_n, n_16084);
  or g47839 (n_16113, n_16084, wc749);
  not gc749 (wc749, rst_n);
  or g47840 (n_20299, wc750, n_17076);
  not gc750 (wc750, \out_fifo[0][0] [4]);
  nand g47841 (n_16115, rst_n, n_16088);
  nand g47842 (n_16118, rst_n, n_16081);
  nand g47843 (n_16523, n_17902, n_22990);
  or g47844 (n_20298, wc751, n_17077);
  not gc751 (wc751, \out_fifo[1][0] [4]);
  or g47845 (n_20297, wc752, n_17079);
  not gc752 (wc752, \out_fifo[5][0] [4]);
  or g47846 (n_20200, wc753, n_17078);
  not gc753 (wc753, \out_fifo[4][1] [0]);
  or g47847 (n_20201, wc754, n_17079);
  not gc754 (wc754, \out_fifo[5][1] [0]);
  or g47848 (n_20202, wc755, n_17077);
  not gc755 (wc755, \out_fifo[1][1] [0]);
  or g47849 (n_20203, wc756, n_17076);
  not gc756 (wc756, \out_fifo[0][1] [0]);
  or g47850 (n_20296, wc757, n_17078);
  not gc757 (wc757, \out_fifo[4][0] [4]);
  nand g47853 (n_16209, n_24564, n_24565);
  or g47854 (n_20205, wc758, n_17068);
  not gc758 (wc758, \out_fifo[7][1] [0]);
  or g47855 (n_20206, wc759, n_17070);
  not gc759 (wc759, \out_fifo[2][1] [0]);
  or g47856 (n_20207, wc760, n_17072);
  not gc760 (wc760, \out_fifo[3][1] [0]);
  or g47857 (n_20208, wc761, n_17074);
  not gc761 (wc761, \out_fifo[6][1] [0]);
  or g47858 (n_16119, n_16081, wc762);
  not gc762 (wc762, rst_n);
  nand g47859 (n_24566, n_16157, n_16166);
  or g47860 (n_24567, n_16157, n_16166);
  nand g47861 (n_16167, n_24566, n_24567);
  nand g47862 (n_16121, rst_n, n_16094);
  or g47863 (n_16122, n_16094, wc763);
  not gc763 (wc763, rst_n);
  nand g47864 (n_16124, rst_n, n_16090);
  or g47865 (n_16125, n_16090, wc764);
  not gc764 (wc764, rst_n);
  nand g47866 (n_16127, rst_n, n_16086);
  or g47867 (n_20248, wc765, n_17078);
  not gc765 (wc765, \out_fifo[4][0] [1]);
  or g47868 (n_20249, wc766, n_17079);
  not gc766 (wc766, \out_fifo[5][0] [1]);
  or g47869 (n_20250, wc767, n_17077);
  not gc767 (wc767, \out_fifo[1][0] [1]);
  or g47870 (n_20251, wc768, n_17076);
  not gc768 (wc768, \out_fifo[0][0] [1]);
  or g47871 (n_16128, n_16086, wc769);
  not gc769 (wc769, rst_n);
  or g47872 (n_20253, wc770, n_17068);
  not gc770 (wc770, \out_fifo[7][0] [1]);
  or g47873 (n_20254, wc771, n_17070);
  not gc771 (wc771, \out_fifo[2][0] [1]);
  or g47874 (n_20255, wc772, n_17072);
  not gc772 (wc772, \out_fifo[3][0] [1]);
  or g47875 (n_20256, wc773, n_17074);
  not gc773 (wc773, \out_fifo[6][0] [1]);
  nand g47876 (n_16130, rst_n, n_16092);
  or g47877 (n_16131, n_16092, wc774);
  not gc774 (wc774, rst_n);
  or g47879 (n_16108, data_parity_mem[1], n_17848);
  nand g47880 (n_23038, n_17384, n_16250);
  nand g47881 (n_16936, n_18813, n_18814);
  or g47882 (n_18903, n_16224, n_16249);
  or g47883 (n_17070, n_17067, n_17069);
  nand g47884 (n_18424, \data_stack_mem[8] [6], n_17043);
  nand g47885 (n_22990, n_17416, n_16483);
  or g47888 (n_16116, out_fifo_write_pointer[2], n_18100);
  nand g47889 (n_18101, out_fifo_write_pointer[2], n_18358);
  nand g47890 (n_24568, n_16504, n_16537);
  or g47891 (n_24569, n_16504, n_16537);
  nand g47892 (n_16538, n_24568, n_24569);
  nand g47894 (n_18301, n_18299, n_18300);
  nand g47896 (n_23008, n_17447, n_16459);
  nand g47897 (n_19470, n_17265, n_16225);
  or g47898 (n_19407, wc775, n_17031);
  not gc775 (wc775, sh_reg_in[3]);
  or g47899 (n_19425, wc776, n_16249);
  not gc776 (wc776, \data_stack_mem[2] [1]);
  nand g47903 (n_16600, n_24570, n_24571);
  nand g47905 (n_18418, \data_stack_mem[8] [5], n_17043);
  nand g47907 (n_24572, n_16206, n_16207);
  or g47908 (n_24573, n_16206, n_16207);
  nand g47909 (n_16208, n_24572, n_24573);
  or g47910 (n_21000, n_20997, wc777);
  not gc777 (wc777, n_16175);
  nand g47911 (n_18412, \data_stack_mem[8] [4], n_17043);
  or g47913 (n_18518, n_16182, wc778);
  not gc778 (wc778, n_18512);
  nand g47916 (n_16278, n_24574, n_24575);
  nand g47917 (n_18406, \data_stack_mem[8] [3], n_17043);
  or g47918 (n_19419, wc779, n_17031);
  not gc779 (wc779, sh_reg_in[4]);
  or g47919 (n_19413, wc780, n_17031);
  not gc780 (wc780, sh_reg_in[1]);
  or g47920 (n_19401, wc781, n_17031);
  not gc781 (wc781, sh_reg_in[2]);
  or g47921 (n_19395, wc782, n_17031);
  not gc782 (wc782, sh_reg_in[0]);
  or g47923 (n_19383, wc783, n_17031);
  not gc783 (wc783, sh_reg_in[7]);
  or g47924 (n_19377, wc784, n_17031);
  not gc784 (wc784, sh_reg_in[6]);
  or g47925 (n_19371, wc785, n_17031);
  not gc785 (wc785, sh_reg_in[5]);
  or g47926 (n_19311, wc786, n_16985);
  not gc786 (wc786, sh_reg_in[7]);
  or g47928 (n_19305, wc787, n_16985);
  not gc787 (wc787, sh_reg_in[6]);
  or g47929 (n_18346, n_16483, n_16437);
  nand g47930 (n_18400, \data_stack_mem[8] [0], n_17043);
  nand g47933 (n_16443, n_24576, n_24577);
  or g47934 (n_19299, wc788, n_16985);
  not gc788 (wc788, sh_reg_in[1]);
  or g47935 (n_23021, data_stack_pointer[4], n_18443);
  or g47936 (n_19293, wc789, n_16985);
  not gc789 (wc789, sh_reg_in[0]);
  nand g47937 (n_18394, \data_stack_mem[8] [2], n_17043);
  or g47940 (n_19281, wc790, n_16985);
  not gc790 (wc790, sh_reg_in[2]);
  or g47941 (n_19275, wc791, n_16985);
  not gc791 (wc791, sh_reg_in[3]);
  or g47942 (n_19269, wc792, n_16985);
  not gc792 (wc792, sh_reg_in[4]);
  or g47943 (n_19263, wc793, n_16985);
  not gc793 (wc793, sh_reg_in[5]);
  nand g47944 (n_16140, n_18387, n_18388);
  or g47946 (n_17074, n_17067, n_17073);
  nand g47949 (n_16365, n_24578, n_24579);
  or g47951 (n_17068, n_17066, n_17067);
  nand g47954 (n_16783, n_24580, n_24581);
  or g47955 (n_17072, n_17067, n_17071);
  or g47956 (n_17964, n_17963, wc794);
  not gc794 (wc794, rst_n);
  or g47957 (n_17848, data_parity_mem[3], n_17847);
  or g47959 (n_19142, data_stack_pointer[3], n_16949);
  or g47960 (n_19135, wc795, n_16949);
  not gc795 (wc795, n_16928);
  or g47961 (n_19132, wc796, n_16949);
  not gc796 (wc796, n_16141);
  or g47964 (n_19461, n_16225, n_16200);
  nand g47966 (n_18568, n_18566, n_18567);
  or g47967 (n_16997, n_17851, n_16949);
  nand g47969 (n_18892, data_parity_mem[2], n_16974);
  or g47971 (n_16088, out_fifo_write_pointer[2], n_18358);
  nand g47972 (n_18886, \data_stack_mem[2] [7], n_16974);
  nand g47974 (n_18880, \data_stack_mem[2] [4], n_16974);
  or g47975 (n_16090, out_fifo_write_pointer[2], n_18361);
  nand g47976 (n_18874, \data_stack_mem[2] [3], n_16974);
  nand g47978 (n_18868, \data_stack_mem[2] [5], n_16974);
  nand g47980 (n_18862, \data_stack_mem[2] [6], n_16974);
  or g47981 (n_18558, data_stack_pointer[0], n_18556);
  nand g47982 (n_18856, \data_stack_mem[2] [1], n_16974);
  nand g47983 (n_23023, data_stack_pointer[4], n_17715);
  nand g47984 (n_18850, \data_stack_mem[2] [0], n_16974);
  nand g47985 (n_24582, n_16159, n_16165);
  or g47986 (n_24583, n_16159, n_16165);
  nand g47987 (n_16166, n_24582, n_24583);
  or g47988 (n_18465, data_stack_pointer[2], n_18464);
  nand g47989 (n_18844, \data_stack_mem[2] [2], n_16974);
  or g47990 (n_17076, n_17069, n_17075);
  nand g47991 (n_18838, data_parity_mem[8], n_17043);
  or g47992 (n_18912, \data_stack_mem[2] [1], wc797);
  not gc797 (wc797, n_17265);
  nand g47993 (n_18832, data_parity_mem[0], n_16930);
  or g47994 (n_17077, n_17071, n_17075);
  or g47996 (n_18323, n_16438, n_16459);
  nand g47998 (n_18826, \data_stack_mem[0] [7], n_16930);
  or g47999 (n_18911, wc798, n_17265);
  not gc798 (wc798, \data_stack_mem[2] [1]);
  or g48000 (n_17079, n_17066, n_17075);
  nand g48001 (n_18820, \data_stack_mem[0] [1], n_16930);
  or g48002 (n_17078, n_17073, n_17075);
  nand g48003 (n_18814, \data_stack_mem[0] [2], n_16930);
  or g48004 (n_18444, data_stack_pointer[3], n_18443);
  nand g48005 (n_18808, \data_stack_mem[0] [3], n_16930);
  or g48006 (n_16092, out_fifo_write_pointer[2], n_17963);
  nand g48007 (n_18802, \data_stack_mem[0] [4], n_16930);
  nand g48008 (n_18313, n_18311, n_18312);
  nand g48009 (n_18796, \data_stack_mem[0] [5], n_16930);
  or g48010 (n_18033, n_18031, n_18032);
  nand g48011 (n_18790, \data_stack_mem[0] [0], n_16930);
  or g48012 (n_16950, n_16141, n_16949);
  nand g48013 (n_18784, \data_stack_mem[0] [6], n_16930);
  or g48014 (n_16094, out_fifo_write_pointer[2], n_18367);
  nand g48015 (n_18436, \data_stack_mem[8] [1], n_17043);
  nand g48017 (n_18430, \data_stack_mem[8] [7], n_17043);
  or g48018 (n_16962, n_16928, n_16949);
  or g48019 (n_18904, n_16200, wc799);
  not gc799 (wc799, n_16249);
  or g48021 (n_17847, data_parity_mem[9], n_17846);
  nand g48022 (n_24584, n_16161, n_16164);
  or g48023 (n_24585, n_16161, n_16164);
  nand g48024 (n_16165, n_24584, n_24585);
  or g48026 (n_17075, out_fifo_read_pointer[1], n_16105);
  or g48027 (n_17067, wc800, n_16105);
  not gc800 (wc800, out_fifo_read_pointer[1]);
  nand g48028 (n_24586, n_16199, n_16205);
  or g48029 (n_24587, n_16199, n_16205);
  nand g48030 (n_16206, n_24586, n_24587);
  nand g48031 (n_24588, n_16501, n_16536);
  or g48032 (n_24589, n_16501, n_16536);
  nand g48033 (n_16537, n_24588, n_24589);
  or g48034 (n_17031, n_16142, n_16984);
  or g48035 (n_16949, wc801, n_16948);
  not gc801 (wc801, data_stack_pointer[0]);
  or g48038 (n_24591, wc802, n_16362);
  not gc802 (wc802, n_16356);
  or g48039 (n_24592, n_16356, wc803);
  not gc803 (wc803, n_16362);
  nand g48040 (n_16363, n_24591, n_24592);
  nand g48046 (n_16599, n_24594, n_24595);
  nand g48050 (n_17944, n_17942, n_17943);
  or g48051 (n_18367, n_16083, out_fifo_write_pointer[0]);
  or g48052 (n_17965, wc804, n_17245);
  not gc804 (wc804, n_17055);
  or g48053 (n_17963, wc805, n_16083);
  not gc805 (wc805, out_fifo_write_pointer[0]);
  or g48054 (n_18100, n_17245, n_17055);
  or g48056 (n_19477, wc806, n_16984);
  not gc806 (wc806, n_16141);
  or g48057 (n_19474, wc807, n_16984);
  not gc807 (wc807, n_16928);
  nand g48058 (n_16483, n_17899, n_22987);
  or g48059 (n_18361, n_16078, out_fifo_write_pointer[0]);
  or g48061 (n_24597, wc808, n_16276);
  not gc808 (wc808, n_16270);
  or g48062 (n_24598, n_16270, wc809);
  not gc809 (wc809, n_16276);
  nand g48063 (n_16277, n_24597, n_24598);
  or g48064 (n_18032, n_18029, n_18030);
  or g48065 (n_16985, n_17373, n_16984);
  or g48066 (n_18031, n_18027, n_18028);
  nand g48071 (n_16782, n_24599, n_24600);
  or g48074 (n_19147, wc810, n_16984);
  not gc810 (wc810, n_16142);
  or g48075 (n_19143, n_16150, n_16948);
  or g48076 (n_19105, data_stack_pointer[0], n_16984);
  nand g48077 (n_17065, n_16105, n_18919);
  nand g48078 (n_17043, n_16133, n_18382);
  nand g48079 (n_17064, n_16105, n_18916);
  or g48080 (n_18387, data_stack_pointer[0], n_16139);
  nand g48081 (n_17063, n_16105, n_18898);
  or g48082 (n_18393, wc811, n_17042);
  not gc811 (wc811, sh_reg_in[2]);
  or g48083 (n_18399, wc812, n_17042);
  not gc812 (wc812, sh_reg_in[0]);
  or g48084 (n_18405, wc813, n_17042);
  not gc813 (wc813, sh_reg_in[3]);
  or g48086 (n_18885, wc814, n_16973);
  not gc814 (wc814, sh_reg_in[7]);
  or g48087 (n_18879, wc815, n_16973);
  not gc815 (wc815, sh_reg_in[4]);
  or g48088 (n_18574, n_16928, n_16984);
  or g48089 (n_18867, wc816, n_16973);
  not gc816 (wc816, sh_reg_in[5]);
  or g48090 (n_18861, wc817, n_16973);
  not gc817 (wc817, sh_reg_in[6]);
  or g48091 (n_18855, wc818, n_16973);
  not gc818 (wc818, sh_reg_in[1]);
  or g48092 (n_18849, wc819, n_16973);
  not gc819 (wc819, sh_reg_in[0]);
  or g48093 (n_18411, wc820, n_17042);
  not gc820 (wc820, sh_reg_in[4]);
  or g48094 (n_18843, wc821, n_16973);
  not gc821 (wc821, sh_reg_in[2]);
  nand g48097 (n_16459, n_17985, n_17986);
  or g48098 (n_18417, wc822, n_17042);
  not gc822 (wc822, sh_reg_in[5]);
  or g48099 (n_18825, wc823, n_16927);
  not gc823 (wc823, sh_reg_in[7]);
  or g48100 (n_18819, wc824, n_16927);
  not gc824 (wc824, sh_reg_in[1]);
  or g48101 (n_18813, wc825, n_16927);
  not gc825 (wc825, sh_reg_in[2]);
  or g48102 (n_18807, wc826, n_16927);
  not gc826 (wc826, sh_reg_in[3]);
  or g48103 (n_18801, wc827, n_16927);
  not gc827 (wc827, sh_reg_in[4]);
  or g48104 (n_18795, wc828, n_16927);
  not gc828 (wc828, sh_reg_in[5]);
  or g48106 (n_18789, wc829, n_16927);
  not gc829 (wc829, sh_reg_in[0]);
  or g48107 (n_18783, wc830, n_16927);
  not gc830 (wc830, sh_reg_in[6]);
  or g48109 (n_18423, wc831, n_17042);
  not gc831 (wc831, sh_reg_in[6]);
  or g48111 (n_18429, wc832, n_17042);
  not gc832 (wc832, sh_reg_in[7]);
  or g48112 (n_18435, wc833, n_17042);
  not gc833 (wc833, sh_reg_in[1]);
  or g48114 (n_18443, n_16151, n_16139);
  nand g48116 (n_18445, data_stack_pointer[3], n_17059);
  or g48118 (n_18358, wc834, n_16078);
  not gc834 (wc834, out_fifo_write_pointer[0]);
  or g48120 (n_17715, n_17059, wc835);
  not gc835 (wc835, n_18448);
  nand g48122 (n_20997, n_16178, n_16176);
  or g48123 (n_18455, data_stack_pointer[1], n_16139);
  or g48124 (n_16182, wc836, n_18205);
  not gc836 (wc836, n_16181);
  nand g48125 (n_18457, n_17718, data_stack_pointer[1]);
  or g48126 (n_18522, n_18519, n_18520);
  nand g48127 (n_18466, n_17719, data_stack_pointer[2]);
  or g48128 (n_24601, wc837, n_16441);
  not gc837 (wc837, n_16435);
  or g48129 (n_24602, n_16435, wc838);
  not gc838 (wc838, n_16441);
  nand g48130 (n_16442, n_24601, n_24602);
  or g48131 (n_18464, n_16150, n_16139);
  nand g48134 (n_16107, n_16105, n_18586);
  nand g48136 (n_16106, n_16105, n_18583);
  or g48139 (n_16930, n_16929, wc839);
  not gc839 (wc839, n_18580);
  or g48140 (n_16974, n_16929, wc840);
  not gc840 (wc840, n_18571);
  or g48141 (n_18577, n_16141, n_16984);
  or g48142 (n_18873, wc841, n_16973);
  not gc841 (wc841, sh_reg_in[3]);
  nand g48148 (n_18481, n_17747, n_17746);
  or g48149 (n_24605, wc842, n_16434);
  not gc842 (wc842, n_16433);
  or g48150 (n_24606, n_16433, wc843);
  not gc843 (wc843, n_16434);
  nand g48151 (n_16435, n_24605, n_24606);
  nand g48152 (n_18079, n_16772, n_16774);
  or g48153 (n_18583, wc844, n_16069);
  not gc844 (wc844, dout_valid);
  or g48154 (n_18586, sh_reg_out_bit_counter[0], n_16069);
  nand g48156 (n_18220, n_17761, n_16147);
  nand g48157 (n_24607, n_16436, n_16440);
  or g48158 (n_24608, n_16436, n_16440);
  nand g48159 (n_16441, n_24607, n_24608);
  or g48160 (n_20684, wc845, n_16069);
  not gc845 (wc845, sh_reg_out[2]);
  nand g48161 (n_18519, n_18513, n_18514);
  nand g48162 (n_18205, n_17756, n_17755);
  nand g48164 (n_18478, n_17745, n_17744);
  or g48167 (n_18311, n_16359, n_16404);
  or g48168 (n_20636, wc846, n_16069);
  not gc846 (wc846, sh_reg_out[1]);
  or g48169 (n_16179, sh_reg_in[1], n_17917);
  nand g48170 (n_18475, n_17743, n_17742);
  nand g48171 (n_18979, n_18975, n_18976);
  nand g48172 (n_18265, n_18263, n_18264);
  nand g48173 (n_18472, n_17737, n_17736);
  or g48174 (n_16176, sh_reg_in[5], n_17923);
  nand g48175 (n_18978, n_18973, n_18974);
  or g48178 (n_20588, wc847, n_16069);
  not gc847 (wc847, sh_reg_out[25]);
  nand g48179 (n_17985, n_17391, n_16404);
  or g48180 (n_20540, wc848, n_16069);
  not gc848 (wc848, sh_reg_out[20]);
  or g48181 (n_20492, wc849, n_16069);
  not gc849 (wc849, sh_reg_out[7]);
  or g48184 (n_18388, wc850, n_16133);
  not gc850 (wc850, data_stack_pointer[0]);
  or g48185 (n_18898, n_18897, n_16069);
  or g48188 (n_17042, n_18379, n_16135);
  nand g48189 (n_18469, n_17735, n_17734);
  or g48192 (n_20444, wc851, n_16069);
  not gc851 (wc851, sh_reg_out[6]);
  or g48193 (n_16973, n_18376, n_16135);
  or g48194 (n_16927, n_16143, n_16135);
  nand g48195 (n_17059, n_18253, n_16133);
  nand g48196 (n_24610, n_16676, n_16780);
  or g48197 (n_24611, n_16676, n_16780);
  nand g48198 (n_16781, n_24610, n_24611);
  nand g48199 (n_18337, n_18335, n_18336);
  nand g48200 (n_18027, n_18019, n_18020);
  or g48201 (n_24612, wc852, n_16778);
  not gc852 (wc852, n_16777);
  or g48202 (n_24613, n_16777, wc853);
  not gc853 (wc853, n_16778);
  nand g48203 (n_16779, n_24612, n_24613);
  nand g48206 (n_16773, n_24614, n_24615);
  nand g48207 (n_18029, n_18023, n_18024);
  or g48208 (n_24616, wc854, n_16269);
  not gc854 (wc854, n_16268);
  or g48209 (n_24617, n_16268, wc855);
  not gc855 (wc855, n_16269);
  nand g48210 (n_16270, n_24616, n_24617);
  nand g48212 (n_24618, n_16271, n_16275);
  or g48213 (n_24619, n_16271, n_16275);
  nand g48214 (n_16276, n_24618, n_24619);
  or g48215 (n_20396, wc856, n_16069);
  not gc856 (wc856, sh_reg_out[5]);
  nand g48216 (n_16929, n_18250, n_16133);
  nand g48218 (n_22987, n_17411, n_16379);
  or g48219 (n_18298, n_16379, n_16358);
  or g48220 (n_19676, wc857, n_16069);
  not gc857 (wc857, sh_reg_out[10]);
  nand g48221 (n_17719, n_16133, n_18091);
  nand g48222 (n_17718, n_16133, n_18088);
  or g48223 (n_16083, out_fifo_write_pointer[1], n_18040);
  or g48224 (n_17057, n_16133, wc858);
  not gc858 (wc858, n_18046);
  or g48225 (n_19724, wc859, n_16069);
  not gc859 (wc859, sh_reg_out[12]);
  or g48226 (n_19772, wc860, n_16069);
  not gc860 (wc860, sh_reg_out[13]);
  or g48227 (n_17055, wc861, n_18040);
  not gc861 (wc861, out_fifo_write_pointer[0]);
  or g48228 (n_19820, wc862, n_16069);
  not gc862 (wc862, sh_reg_out[14]);
  or g48229 (n_19868, wc863, n_16069);
  not gc863 (wc863, sh_reg_out[11]);
  nand g48230 (n_17943, out_fifo_read_pointer[2], n_17290);
  or g48231 (n_17942, n_17071, n_17290);
  or g48232 (n_19916, wc864, n_16069);
  not gc864 (wc864, sh_reg_out[16]);
  nand g48233 (n_24620, out_fifo_read_pointer[1], n_17300);
  or g48234 (n_24621, out_fifo_read_pointer[1], n_17300);
  nand g48235 (n_17732, n_24620, n_24621);
  nand g48246 (n_18526, n_17759, n_17758);
  or g48247 (n_20348, wc865, n_16069);
  not gc865 (wc865, sh_reg_out[4]);
  nand g48248 (n_18241, n_17762, n_16352);
  or g48249 (n_19964, wc866, n_16069);
  not gc866 (wc866, sh_reg_out[17]);
  nand g48252 (n_24628, n_16593, n_16597);
  or g48253 (n_24629, n_16593, n_16597);
  nand g48254 (n_16598, n_24628, n_24629);
  or g48255 (n_20012, wc867, n_16069);
  not gc867 (wc867, sh_reg_out[27]);
  nand g48256 (n_24630, n_16357, n_16361);
  or g48257 (n_24631, n_16357, n_16361);
  nand g48258 (n_16362, n_24630, n_24631);
  nand g48259 (n_24632, out_fifo_write_pointer[0], n_18040);
  or g48260 (n_24633, out_fifo_write_pointer[0], n_18040);
  nand g48261 (n_17724, n_24632, n_24633);
  or g48262 (n_24634, wc868, n_16591);
  not gc868 (wc868, n_16590);
  or g48263 (n_24635, n_16590, wc869);
  not gc869 (wc869, n_16591);
  nand g48264 (n_16592, n_24634, n_24635);
  nand g48265 (n_17723, n_17970, n_17971);
  nand g48268 (n_16946, n_24636, n_24637);
  or g48269 (n_16948, n_16135, n_16137);
  or g48270 (n_20060, wc870, n_16069);
  not gc870 (wc870, sh_reg_out[28]);
  or g48271 (n_16984, n_18370, n_16135);
  or g48272 (n_24638, wc871, n_16353);
  not gc871 (wc871, n_16352);
  or g48273 (n_24639, n_16352, wc872);
  not gc872 (wc872, n_16353);
  nand g48274 (n_16354, n_24638, n_24639);
  or g48275 (n_20108, wc873, n_16069);
  not gc873 (wc873, sh_reg_out[15]);
  or g48276 (n_20156, wc874, n_16069);
  not gc874 (wc874, sh_reg_out[19]);
  nand g48277 (n_24640, n_16200, n_16204);
  or g48278 (n_24641, n_16200, n_16204);
  nand g48279 (n_16205, n_24640, n_24641);
  or g48280 (n_16183, sh_reg_in[0], n_16178);
  or g48281 (n_16105, wc875, n_17286);
  not gc875 (wc875, n_17716);
  or g48282 (n_24642, wc876, n_16535);
  not gc876 (wc876, n_16503);
  or g48283 (n_24643, n_16503, wc877);
  not gc877 (wc877, n_16535);
  nand g48284 (n_16536, n_24642, n_24643);
  nand g48285 (n_18277, n_18275, n_18276);
  nand g48286 (n_17390, n_16143, n_16898);
  or g48287 (n_17846, data_parity_mem[0], n_17845);
  or g48288 (n_20300, wc878, n_16069);
  not gc878 (wc878, sh_reg_out[3]);
  nand g48289 (n_16164, n_18354, n_18355);
  or g48291 (n_20204, wc879, n_16069);
  not gc879 (wc879, sh_reg_out[9]);
  nand g48292 (n_18289, n_18287, n_18288);
  or g48295 (n_20252, wc880, n_16069);
  not gc880 (wc880, sh_reg_out[0]);
  or g48296 (n_17845, data_parity_mem[5], n_17844);
  nand g48297 (n_19068, n_19064, n_19065);
  or g48298 (n_19066, \data_stack_mem[4] [7], wc881);
  not gc881 (wc881, n_16156);
  nand g48299 (n_17747, n_16682, n_18154);
  or g48300 (n_18287, n_16273, n_16319);
  or g48302 (n_24645, wc882, n_16197);
  not gc882 (wc882, n_16196);
  or g48303 (n_24646, n_16196, wc883);
  not gc883 (wc883, n_16197);
  nand g48304 (n_16198, n_24645, n_24646);
  nand g48305 (n_18142, n_17741, n_16196);
  or g48306 (n_19063, \data_stack_mem[8] [7], wc884);
  not gc884 (wc884, n_16146);
  or g48307 (n_18448, data_stack_pointer[3], n_16924);
  or g48308 (n_18976, \data_stack_mem[4] [1], wc885);
  not gc885 (wc885, n_16156);
  nand g48309 (n_16275, n_16273, n_16274);
  nand g48310 (n_17737, n_17890, n_16203);
  or g48311 (n_18088, data_stack_pointer[0], n_16924);
  nand g48312 (n_18354, n_17635, \data_stack_mem[0] [0]);
  nand g48313 (n_16361, n_16359, n_16360);
  or g48314 (n_18973, \data_stack_mem[8] [1], wc886);
  not gc886 (wc886, n_16146);
  or g48316 (n_18091, wc887, n_16924);
  not gc887 (wc887, n_16150);
  nand g48317 (n_16379, n_17896, n_22984);
  nand g48320 (n_16945, n_24647, n_24648);
  or g48321 (n_24649, wc888, n_16266);
  not gc888 (wc888, n_16265);
  or g48322 (n_24650, n_16265, wc889);
  not gc889 (wc889, n_16266);
  nand g48323 (n_16267, n_24649, n_24650);
  nand g48324 (n_18945, n_18941, n_18942);
  nand g48325 (n_16404, n_17949, n_17950);
  or g48326 (n_18943, \data_stack_mem[4] [6], wc890);
  not gc890 (wc890, n_16156);
  nand g48327 (n_17735, n_16596, n_18106);
  or g48328 (n_24651, wc891, n_16431);
  not gc891 (wc891, n_16430);
  or g48329 (n_24652, n_16430, wc892);
  not gc892 (wc892, n_16431);
  nand g48330 (n_16432, n_24651, n_24652);
  or g48331 (n_18940, \data_stack_mem[8] [6], wc893);
  not gc893 (wc893, n_16146);
  nand g48332 (n_17729, n_17859, n_17860);
  nand g48333 (n_18121, n_17740, n_16587);
  or g48334 (n_18040, wc894, n_16077);
  not gc894 (wc894, sh_reg_in[8]);
  or g48335 (n_24653, wc895, n_16775);
  not gc895 (wc895, n_16774);
  or g48336 (n_24654, n_16774, wc896);
  not gc896 (wc896, n_16775);
  nand g48337 (n_16776, n_24653, n_24654);
  nand g48338 (n_16440, n_16438, n_16439);
  nand g48339 (n_16780, n_16681, n_16682);
  or g48340 (n_18336, wc897, n_16202);
  not gc897 (wc897, n_16163);
  or g48341 (n_18335, n_18355, n_16201);
  or g48342 (n_23002, sh_reg_in[4], n_17922);
  or g48344 (n_18020, \data_stack_mem[8] [5], wc898);
  not gc898 (wc898, n_16146);
  or g48345 (n_18264, wc899, n_16202);
  not gc899 (wc899, n_16180);
  or g48346 (n_18253, wc900, n_16924);
  not gc900 (wc900, n_16151);
  nand g48347 (n_18028, n_18021, n_18022);
  nand g48348 (n_19038, n_19034, n_19035);
  or g48349 (n_19036, \data_stack_mem[4] [2], wc901);
  not gc901 (wc901, n_16156);
  nand g48350 (n_17743, n_17950, n_16274);
  or g48351 (n_16135, n_16077, n_16134);
  or g48352 (n_19033, \data_stack_mem[8] [2], wc902);
  not gc902 (wc902, n_16146);
  or g48353 (n_18276, n_16273, wc903);
  not gc903 (wc903, n_16293);
  or g48356 (n_18024, \data_stack_mem[4] [5], wc904);
  not gc904 (wc904, n_16156);
  nand g48357 (n_18196, n_17754, n_16265);
  nand g48358 (n_16204, n_16202, n_16203);
  nand g48359 (n_24655, out_fifo_read_pointer[0], n_16103);
  or g48360 (n_24656, out_fifo_read_pointer[0], n_16103);
  nand g48361 (n_17731, n_24655, n_24656);
  nand g48362 (n_19008, n_19004, n_19005);
  nand g48363 (n_16535, n_16522, n_18043);
  or g48364 (n_19006, \data_stack_mem[4] [4], wc905);
  not gc905 (wc905, n_16156);
  nand g48365 (n_17745, n_16439, n_18151);
  nand g48366 (n_18030, n_18025, n_18026);
  or g48367 (n_19003, \data_stack_mem[8] [4], wc906);
  not gc906 (wc906, n_16146);
  nand g48368 (n_16133, n_16077, rst_n);
  or g48369 (n_24657, wc907, n_16588);
  not gc907 (wc907, n_16587);
  or g48370 (n_24658, n_16587, wc908);
  not gc908 (wc908, n_16588);
  nand g48371 (n_16589, n_24657, n_24658);
  nand g48372 (n_18175, n_17753, n_16430);
  nand g48373 (n_18060, n_16501, n_18059);
  or g48374 (n_18517, \data_stack_mem[4] [0], wc909);
  not gc909 (wc909, n_16156);
  or g48375 (n_17286, n_16068, wc910);
  not gc910 (wc910, rst_n);
  nand g48376 (n_17756, n_16180, n_17977);
  nand g48377 (n_16069, n_16068, rst_n);
  nand g48378 (n_16597, n_16595, n_16596);
  or g48379 (n_18513, \data_stack_mem[8] [0], wc911);
  not gc911 (wc911, n_16146);
  nand g48380 (n_17970, n_17722, n_16100);
  nand g48381 (n_19098, n_19094, n_19095);
  or g48382 (n_19096, \data_stack_mem[4] [3], wc912);
  not gc912 (wc912, n_16156);
  nand g48383 (n_18520, n_18515, n_18516);
  nand g48384 (n_17759, n_17986, n_16360);
  nand g48385 (n_16898, n_17763, n_16143);
  or g48386 (n_19093, \data_stack_mem[8] [3], wc913);
  not gc913 (wc913, n_16146);
  nand g48389 (n_16944, n_24659, n_24660);
  or g48390 (n_16203, wc914, n_16162);
  not gc914 (wc914, \data_stack_mem[0] [1]);
  nand g48391 (n_18897, sh_reg_out_bit_counter[4], n_16067);
  or g48392 (n_18286, wc915, n_16272);
  not gc915 (wc915, n_16319);
  or g48393 (n_18379, n_17387, wc916);
  not gc916 (wc916, n_16136);
  or g48394 (n_19095, \data_stack_mem[5] [3], wc917);
  not gc917 (wc917, n_16154);
  or g48395 (n_19094, \data_stack_mem[6] [3], wc918);
  not gc918 (wc918, n_16152);
  nand g48396 (n_16359, n_16162, n_16358);
  or g48397 (n_16360, wc919, n_16162);
  not gc919 (wc919, \data_stack_mem[0] [3]);
  nand g48398 (n_22984, n_17442, n_16293);
  nand g48399 (n_18059, n_16162, n_17303);
  nand g48400 (n_18046, sh_bit_cnt[3], n_16076);
  or g48401 (n_16391, \data_stack_mem[9] [3], wc920);
  not gc920 (wc920, n_16145);
  nand g48402 (n_17727, n_16067, n_17974);
  nand g48403 (n_17949, n_17417, n_16319);
  or g48404 (n_18026, \data_stack_mem[1] [5], wc921);
  not gc921 (wc921, n_16162);
  or g48405 (n_16306, \data_stack_mem[9] [2], wc922);
  not gc922 (wc922, n_16145);
  or g48406 (n_18025, \data_stack_mem[2] [5], wc923);
  not gc923 (wc923, n_16160);
  or g48407 (n_18023, \data_stack_mem[5] [5], wc924);
  not gc924 (wc924, n_16154);
  or g48408 (n_18021, \data_stack_mem[6] [5], wc925);
  not gc925 (wc925, n_16152);
  or g48409 (n_17859, n_17053, n_17858);
  nand g48410 (n_16438, n_16162, n_16437);
  or g48411 (n_16439, wc926, n_16162);
  not gc926 (wc926, \data_stack_mem[0] [4]);
  nand g48412 (n_16202, n_16162, n_16201);
  nand g48413 (n_17722, n_17932, n_16076);
  or g48415 (n_18160, \data_stack_mem[9] [5], wc927);
  not gc927 (wc927, n_16145);
  or g48416 (n_17763, n_17872, n_16173);
  or g48417 (n_16471, \data_stack_mem[9] [4], wc928);
  not gc928 (wc928, n_16145);
  or g48418 (n_18942, \data_stack_mem[5] [6], wc929);
  not gc929 (wc929, n_16154);
  or g48419 (n_18941, \data_stack_mem[6] [6], wc930);
  not gc930 (wc930, n_16152);
  or g48420 (n_17844, data_parity_mem[4], n_17843);
  or g48421 (n_18274, n_16293, n_16272);
  or g48422 (n_18974, \data_stack_mem[6] [1], wc931);
  not gc931 (wc931, n_16152);
  or g48423 (n_16522, wc932, n_16521);
  not gc932 (wc932, n_16162);
  or g48424 (n_18539, wc933, n_16162);
  not gc933 (wc933, \data_stack_mem[0] [5]);
  or g48425 (n_18043, \data_stack_mem[0] [5], n_16162);
  or g48426 (n_16924, wc934, n_16134);
  not gc934 (wc934, n_17296);
  or g48427 (n_18975, \data_stack_mem[5] [1], wc935);
  not gc935 (wc935, n_16154);
  or g48428 (n_16235, \data_stack_mem[9] [1], wc936);
  not gc936 (wc936, n_16145);
  or g48429 (n_16146, n_16145, wc937);
  not gc937 (wc937, n_17953);
  or g48430 (n_19065, \data_stack_mem[5] [7], wc938);
  not gc938 (wc938, n_16154);
  nand g48431 (n_16595, n_16162, n_16594);
  or g48432 (n_16596, wc939, n_16162);
  not gc939 (wc939, \data_stack_mem[0] [6]);
  or g48433 (n_19064, \data_stack_mem[6] [7], wc940);
  not gc940 (wc940, n_16152);
  nand g48434 (n_17761, n_16162, n_17980);
  or g48435 (n_16156, data_stack_pointer[4], wc941);
  not gc941 (wc941, n_17956);
  or g48436 (n_16628, \data_stack_mem[9] [6], wc942);
  not gc942 (wc942, n_16145);
  or g48437 (n_16682, wc943, n_16162);
  not gc943 (wc943, \data_stack_mem[0] [7]);
  or g48438 (n_18516, \data_stack_mem[5] [0], wc944);
  not gc944 (wc944, n_16154);
  or g48439 (n_18515, \data_stack_mem[6] [0], wc945);
  not gc945 (wc945, n_16152);
  nand g48440 (n_16681, n_16162, n_16680);
  or g48441 (n_18355, wc946, n_16163);
  not gc946 (wc946, n_16162);
  or g48442 (n_18514, \data_stack_mem[9] [0], wc947);
  not gc947 (wc947, n_16145);
  or g48443 (n_16274, wc948, n_16162);
  not gc948 (wc948, \data_stack_mem[0] [2]);
  nand g48444 (n_16273, n_16162, n_16272);
  or g48445 (n_17977, wc949, n_16162);
  not gc949 (wc949, \data_stack_mem[0] [0]);
  or g48446 (n_17916, n_16177, n_16173);
  nand g48448 (n_17467, n_16162, n_18037);
  or g48449 (n_16785, \data_stack_mem[9] [7], wc950);
  not gc950 (wc950, n_16145);
  or g48450 (n_17922, n_16174, n_16173);
  or g48451 (n_19034, \data_stack_mem[6] [2], wc951);
  not gc951 (wc951, n_16152);
  or g48452 (n_19035, \data_stack_mem[5] [2], wc952);
  not gc952 (wc952, n_16154);
  or g48454 (n_19005, \data_stack_mem[5] [4], wc953);
  not gc953 (wc953, n_16154);
  or g48455 (n_19004, \data_stack_mem[6] [4], wc954);
  not gc954 (wc954, n_16152);
  or g48456 (n_18262, n_16180, n_16201);
  or g48457 (n_16173, sh_reg_in[3], n_17824);
  or g48458 (n_17799, n_17805, n_17806);
  or g48459 (n_17296, n_16136, n_16926);
  nand g48460 (n_17956, n_16142, n_17298);
  or g48461 (n_16154, data_stack_pointer[4], wc955);
  not gc955 (wc955, n_17926);
  or g48462 (n_16145, data_stack_pointer[4], wc956);
  not gc956 (wc956, n_17929);
  nand g48463 (n_16293, n_17883, n_17884);
  or g48464 (n_17843, data_parity_mem[2], n_17842);
  or g48465 (n_16143, n_16926, n_16141);
  nand g48466 (n_17872, n_17870, n_17871);
  or g48467 (n_17818, sh_reg_out_bit_counter[4], n_17817);
  or g48468 (n_17858, sh_bit_cnt[1], wc957);
  not gc957 (wc957, n_16100);
  or g48469 (n_18022, \data_stack_mem[3] [5], wc958);
  not gc958 (wc958, n_16158);
  or g48470 (n_16099, n_17772, wc959);
  not gc959 (wc959, rst_n);
  nand g48471 (n_17728, n_16066, n_17935);
  nand g48472 (n_17974, sh_reg_out_bit_counter[3], n_16066);
  or g48474 (n_18376, n_16926, n_16928);
  nand g48475 (n_16319, n_17889, n_17890);
  or g48476 (n_16076, sh_bit_cnt[1], n_17893);
  nand g48479 (n_16943, n_24661, n_24662);
  nand g48482 (n_16942, n_24663, n_24664);
  nand g48483 (n_16594, n_17443, n_17908);
  nand g48486 (n_16940, n_24665, n_24666);
  or g48487 (n_17260, \data_stack_mem[7] [3], wc960);
  not gc960 (wc960, n_16148);
  nand g48488 (n_16358, n_17411, n_17899);
  nand g48489 (n_17805, n_17801, n_17802);
  or g48490 (n_16100, sh_bit_cnt[2], sh_bit_cnt[3]);
  nand g48491 (n_17971, sh_bit_cnt[2], n_17053);
  or g48492 (n_16302, \data_stack_mem[7] [2], wc961);
  not gc961 (wc961, n_16148);
  nand g48493 (n_17929, n_17720, data_stack_pointer[3]);
  nand g48494 (n_16201, n_17353, n_17884);
  or g48495 (n_18019, \data_stack_mem[7] [5], wc962);
  not gc962 (wc962, n_16148);
  nand g48496 (n_17860, sh_bit_cnt[1], n_17053);
  or g48497 (n_18972, \data_stack_mem[7] [1], wc963);
  not gc963 (wc963, n_16148);
  or g48498 (n_18512, \data_stack_mem[7] [0], wc964);
  not gc964 (wc964, n_16148);
  nand g48499 (n_17806, n_17803, n_17804);
  nand g48501 (n_17870, n_16174, n_16177);
  or g48502 (n_17824, sh_reg_in[2], n_17823);
  nand g48503 (n_17730, n_16065, n_17863);
  nand g48504 (n_17883, n_16163, n_17353);
  nand g48505 (n_16521, n_17425, n_17905);
  or g48506 (n_17842, data_parity_mem[8], n_17841);
  or g48507 (n_18567, wc965, n_16134);
  not gc965 (wc965, data_stack_pointer[4]);
  nand g48508 (n_17772, n_17053, n_17771);
  nand g48509 (n_16437, n_17416, n_17902);
  nand g48510 (n_17714, n_16928, n_17851);
  nand g48511 (n_17935, sh_reg_out_bit_counter[2], n_16065);
  or g48512 (n_17893, sh_bit_cnt[2], n_17053);
  nand g48513 (n_16272, n_17442, n_17896);
  or g48514 (n_18571, data_stack_pointer[1], n_16134);
  or g48515 (n_16690, \data_stack_mem[7] [7], wc966);
  not gc966 (wc966, n_16148);
  nand g48516 (n_16680, n_17294, n_17911);
  or g48517 (n_17817, sh_reg_out_bit_counter[3], n_17816);
  or g48518 (n_16467, \data_stack_mem[7] [4], wc967);
  not gc967 (wc967, n_16148);
  or g48519 (n_16624, \data_stack_mem[7] [6], wc968);
  not gc968 (wc968, n_16148);
  or g48520 (n_17706, data_stack_pointer[0], n_16136);
  nand g48521 (n_17926, n_16141, n_17298);
  or g48522 (n_17889, n_16180, wc969);
  not gc969 (wc969, n_17369);
  nand g48525 (n_16941, n_24667, n_24668);
  or g48526 (n_18370, wc970, data_stack_pointer[4]);
  not gc970 (wc970, data_stack_pointer[2]);
  nand g48527 (n_17066, out_fifo_read_pointer[2],
       out_fifo_read_pointer[0]);
  or g48528 (n_17801, out_fifo_read_pointer[1], wc971);
  not gc971 (wc971, out_fifo_write_pointer[1]);
  or g48529 (n_17802, wc972, out_fifo_write_pointer[1]);
  not gc972 (wc972, out_fifo_read_pointer[1]);
  or g48530 (n_17803, out_fifo_read_pointer[2], wc973);
  not gc973 (wc973, out_fifo_write_pointer[2]);
  or g48531 (n_17804, wc974, out_fifo_write_pointer[2]);
  not gc974 (wc974, out_fifo_read_pointer[2]);
  nand g48534 (n_16939, n_24669, n_24670);
  or g48535 (n_17884, wc975, \data_stack_mem[1] [1]);
  not gc975 (wc975, \data_stack_mem[0] [1]);
  or g48536 (n_17980, \data_stack_mem[0] [0], \data_stack_mem[1] [0]);
  or g48537 (n_18037, \data_stack_mem[0] [7], \data_stack_mem[1] [7]);
  nand g48538 (n_18154, \data_stack_mem[0] [7], \data_stack_mem[1] [7]);
  or g48539 (n_17823, sh_reg_in[6], sh_reg_in[7]);
  nand g48542 (n_17800, n_24671, n_24672);
  or g48543 (n_17896, wc976, \data_stack_mem[1] [2]);
  not gc976 (wc976, \data_stack_mem[0] [2]);
  or g48544 (n_17069, out_fifo_read_pointer[2],
       out_fifo_read_pointer[0]);
  or g48545 (n_17071, wc977, out_fifo_read_pointer[2]);
  not gc977 (wc977, out_fifo_read_pointer[0]);
  or g48546 (n_17073, out_fifo_read_pointer[0], wc978);
  not gc978 (wc978, out_fifo_read_pointer[2]);
  nand g48547 (n_17245, rst_n, out_fifo_write_pointer[1]);
  nand g48548 (n_18106, \data_stack_mem[0] [6], \data_stack_mem[1] [6]);
  or g48549 (n_17911, \data_stack_mem[0] [7], wc979);
  not gc979 (wc979, \data_stack_mem[1] [7]);
  nand g48550 (n_18547, \data_stack_mem[0] [5], \data_stack_mem[1] [5]);
  or g48551 (n_17908, wc980, \data_stack_mem[1] [6]);
  not gc980 (wc980, \data_stack_mem[0] [6]);
  nand g48552 (n_17953, data_stack_pointer[0], data_stack_pointer[3]);
  nand g48553 (n_18151, \data_stack_mem[0] [4], \data_stack_mem[1] [4]);
  nand g48554 (n_17871, sh_reg_in[4], sh_reg_in[5]);
  or g48555 (n_17841, data_parity_mem[6], data_parity_mem[7]);
  or g48556 (n_17905, wc981, \data_stack_mem[1] [5]);
  not gc981 (wc981, \data_stack_mem[0] [5]);
  nand g48557 (n_16136, data_stack_pointer[3], data_stack_pointer[1]);
  or g48558 (n_16134, sh_reg_in[8], wc982);
  not gc982 (wc982, rst_n);
  or g48559 (n_17816, sh_reg_out_bit_counter[1],
       sh_reg_out_bit_counter[2]);
  nand g48560 (n_17986, \data_stack_mem[0] [3], \data_stack_mem[1] [3]);
  nand g48561 (n_17932, sh_bit_cnt[1], sh_bit_cnt[2]);
  nand g48563 (n_17863, sh_reg_out_bit_counter[0],
       sh_reg_out_bit_counter[1]);
  nand g48564 (n_17771, sh_bit_cnt[0], enable_n);
  or g48565 (n_17851, data_stack_pointer[1], wc983);
  not gc983 (wc983, data_stack_pointer[3]);
  or g48566 (n_17902, wc984, \data_stack_mem[1] [4]);
  not gc984 (wc984, \data_stack_mem[0] [4]);
  nand g48567 (n_17950, \data_stack_mem[0] [2], \data_stack_mem[1] [2]);
  or g48568 (n_17899, wc985, \data_stack_mem[1] [3]);
  not gc985 (wc985, \data_stack_mem[0] [3]);
  nand g48569 (n_17890, \data_stack_mem[0] [1], \data_stack_mem[1] [1]);
  and g48574 (n_24624, n_17729, rst_n);
  and g48579 (n_24590, n_17723, rst_n);
  and g48580 (n_24622, n_17731, rst_n);
  and g48581 (n_24593, n_17724, rst_n);
  and g48582 (n_24596, n_17732, rst_n);
  and g48583 (n_24561, n_17733, rst_n);
  or g48587 (n_16828, wc986, n_16827);
  not gc986 (wc986, n_17354);
  or g48589 (n_24671, wc987, out_fifo_read_pointer[0]);
  not gc987 (wc987, out_fifo_write_pointer[0]);
  or g48590 (n_24672, out_fifo_write_pointer[0], wc988);
  not gc988 (wc988, out_fifo_read_pointer[0]);
  or g48591 (n_24669, wc989, sh_reg_in[1]);
  not gc989 (wc989, sh_reg_in[3]);
  or g48592 (n_24670, sh_reg_in[3], wc990);
  not gc990 (wc990, sh_reg_in[1]);
  or g48593 (n_24667, wc991, sh_reg_in[7]);
  not gc991 (wc991, din);
  or g48594 (n_24668, din, wc992);
  not gc992 (wc992, sh_reg_in[7]);
  or g48595 (n_18557, n_16134, wc993);
  not gc993 (wc993, n_16137);
  or g48596 (n_24665, wc994, sh_reg_in[4]);
  not gc994 (wc994, n_16939);
  or g48597 (n_24666, n_16939, wc995);
  not gc995 (wc995, sh_reg_in[4]);
  or g48598 (n_24663, wc996, sh_reg_in[5]);
  not gc996 (wc996, n_16941);
  or g48599 (n_24664, n_16941, wc997);
  not gc997 (wc997, sh_reg_in[5]);
  or g48600 (n_18250, n_16134, wc998);
  not gc998 (wc998, n_16926);
  or g48601 (n_18263, n_18262, wc999);
  not gc999 (wc999, n_16162);
  or g48602 (n_23013, n_18154, wc1000);
  not gc1000 (wc1000, n_16162);
  or g48603 (n_16103, n_17818, wc1001);
  not gc1001 (wc1001, sh_reg_out_bit_counter[0]);
  or g48604 (n_18275, n_18274, wc1002);
  not gc1002 (wc1002, n_16162);
  or g48605 (n_18288, n_18286, wc1003);
  not gc1003 (wc1003, n_16162);
  or g48606 (n_17923, n_17922, wc1004);
  not gc1004 (wc1004, sh_reg_in[4]);
  or g48607 (n_16178, n_17916, wc1005);
  not gc1005 (wc1005, sh_reg_in[1]);
  or g48608 (n_17917, n_17916, wc1006);
  not gc1006 (wc1006, sh_reg_in[0]);
  or g48609 (n_24661, wc1007, sh_reg_in[2]);
  not gc1007 (wc1007, n_16942);
  or g48610 (n_24662, n_16942, wc1008);
  not gc1008 (wc1008, sh_reg_in[2]);
  or g48611 (n_16078, n_18040, wc1009);
  not gc1009 (wc1009, out_fifo_write_pointer[1]);
  or g48612 (n_18300, n_16359, wc1010);
  not gc1010 (wc1010, n_16379);
  or g48613 (n_18310, n_16358, wc1011);
  not gc1011 (wc1011, n_16404);
  or g48614 (n_16175, n_23002, wc1012);
  not gc1012 (wc1012, sh_reg_in[5]);
  or g48615 (n_18197, n_18196, wc1013);
  not gc1013 (wc1013, n_16266);
  or g48616 (n_18176, n_18175, wc1014);
  not gc1014 (wc1014, n_16431);
  or g48617 (n_24614, wc1015, n_16667);
  not gc1015 (wc1015, n_16772);
  or g48618 (n_24615, n_16772, wc1016);
  not gc1016 (wc1016, n_16667);
  or g48619 (n_18143, n_18142, wc1017);
  not gc1017 (wc1017, n_16197);
  or g48620 (n_18122, n_18121, wc1018);
  not gc1018 (wc1018, n_16588);
  or g48621 (n_18061, n_18060, wc1019);
  not gc1019 (wc1019, n_16502);
  or g48622 (n_16139, wc1020, n_16135);
  not gc1020 (wc1020, n_17296);
  or g48623 (n_18382, n_16135, wc1021);
  not gc1021 (wc1021, n_17387);
  or g48624 (n_18580, wc1022, n_16135);
  not gc1022 (wc1022, n_17714);
  or g48625 (n_18919, wc1023, n_16069);
  not gc1023 (wc1023, n_17728);
  or g48626 (n_18916, wc1024, n_16069);
  not gc1024 (wc1024, n_17727);
  and g48627 (n_24603, wc1025, sh_reg_out[24]);
  not gc1025 (wc1025, n_16069);
  and g48628 (n_24604, wc1026, sh_reg_out[26]);
  not gc1026 (wc1026, n_16069);
  and g48629 (n_24609, wc1027, sh_reg_out[23]);
  not gc1027 (wc1027, n_16069);
  and g48630 (n_24623, n_17730, wc1028);
  not gc1028 (wc1028, n_16069);
  and g48631 (n_24625, wc1029, sh_reg_out[8]);
  not gc1029 (wc1029, n_16069);
  and g48632 (n_24626, wc1030, sh_reg_out[18]);
  not gc1030 (wc1030, n_16069);
  and g48633 (n_24627, wc1031, sh_reg_out[21]);
  not gc1031 (wc1031, n_16069);
  and g48634 (n_24644, wc1032, sh_reg_out[22]);
  not gc1032 (wc1032, n_16069);
  or g48635 (n_16225, wc1033, n_18337);
  not gc1033 (wc1033, n_16203);
  or g48636 (n_16294, wc1034, n_18277);
  not gc1034 (wc1034, n_16274);
  or g48637 (n_18299, n_18298, wc1035);
  not gc1035 (wc1035, n_16162);
  or g48638 (n_16250, wc1036, n_18265);
  not gc1036 (wc1036, n_16203);
  or g48639 (n_16320, wc1037, n_18289);
  not gc1037 (wc1037, n_16274);
  or g48640 (n_18312, n_18310, wc1038);
  not gc1038 (wc1038, n_16162);
  or g48641 (n_16332, n_18475, wc1039);
  not gc1039 (wc1039, n_16296);
  or g48642 (n_18198, n_18197, wc1040);
  not gc1040 (wc1040, n_16269);
  or g48643 (n_16495, n_18478, wc1041);
  not gc1041 (wc1041, n_16458);
  or g48644 (n_18177, n_18176, wc1042);
  not gc1042 (wc1042, n_16433);
  or g48645 (n_18221, n_18220, wc1043);
  not gc1043 (wc1043, n_16153);
  or g48646 (n_16787, n_18481, wc1044);
  not gc1044 (wc1044, n_16677);
  or g48647 (n_18080, n_18079, wc1045);
  not gc1045 (wc1045, n_16775);
  or g48648 (n_16259, n_18472, wc1046);
  not gc1046 (wc1046, n_16224);
  or g48649 (n_18144, n_18143, wc1047);
  not gc1047 (wc1047, n_16199);
  or g48650 (n_16654, n_18469, wc1048);
  not gc1048 (wc1048, n_16616);
  or g48651 (n_18123, n_18122, wc1049);
  not gc1049 (wc1049, n_16590);
  or g48652 (n_18062, n_18061, wc1050);
  not gc1050 (wc1050, n_16503);
  or g48653 (n_16417, n_18526, wc1051);
  not gc1051 (wc1051, n_16382);
  or g48654 (n_18242, n_18241, wc1052);
  not gc1052 (wc1052, n_16355);
  or g48655 (n_18566, wc1053, n_16948);
  not gc1053 (wc1053, n_17706);
  or g48656 (n_18556, wc1054, n_16948);
  not gc1054 (wc1054, n_16136);
  or g48657 (n_24659, wc1055, sh_reg_in[6]);
  not gc1055 (wc1055, n_16943);
  or g48658 (n_24660, n_16943, wc1056);
  not gc1056 (wc1056, sh_reg_in[6]);
  or g48659 (n_19150, n_16984, wc1057);
  not gc1057 (wc1057, n_17373);
  or g48660 (n_16079, n_18358, wc1058);
  not gc1058 (wc1058, out_fifo_write_pointer[2]);
  or g48661 (n_16081, n_18361, wc1059);
  not gc1059 (wc1059, out_fifo_write_pointer[2]);
  or g48662 (n_16084, n_17963, wc1060);
  not gc1060 (wc1060, out_fifo_write_pointer[2]);
  or g48663 (n_16086, n_18367, wc1061);
  not gc1061 (wc1061, out_fifo_write_pointer[2]);
  or g48664 (n_18348, n_16438, wc1062);
  not gc1062 (wc1062, n_16483);
  or g48665 (n_18322, n_16437, wc1063);
  not gc1063 (wc1063, n_16459);
  or g48666 (n_19037, n_16332, wc1064);
  not gc1064 (wc1064, n_19033);
  or g48667 (n_18199, n_18198, wc1065);
  not gc1065 (wc1065, n_16271);
  or g48668 (n_19007, n_16495, wc1066);
  not gc1066 (wc1066, n_19003);
  or g48669 (n_18178, n_18177, wc1067);
  not gc1067 (wc1067, n_16434);
  or g48670 (n_18222, n_18221, wc1068);
  not gc1068 (wc1068, n_16155);
  or g48671 (n_24599, wc1069, n_16781);
  not gc1069 (wc1069, n_16779);
  or g48672 (n_24600, n_16779, wc1070);
  not gc1070 (wc1070, n_16781);
  or g48673 (n_19067, n_16787, wc1071);
  not gc1071 (wc1071, n_19063);
  or g48674 (n_18081, n_18080, wc1072);
  not gc1072 (wc1072, n_16777);
  or g48675 (n_18977, n_16259, wc1073);
  not gc1073 (wc1073, n_18972);
  or g48676 (n_18145, n_18144, wc1074);
  not gc1074 (wc1074, n_16207);
  or g48677 (n_24594, wc1075, n_16598);
  not gc1075 (wc1075, n_16592);
  or g48678 (n_24595, n_16592, wc1076);
  not gc1076 (wc1076, n_16598);
  or g48679 (n_18944, n_16654, wc1077);
  not gc1077 (wc1077, n_18940);
  or g48680 (n_18124, n_18123, wc1078);
  not gc1078 (wc1078, n_16591);
  or g48681 (n_18063, n_18062, wc1079);
  not gc1079 (wc1079, n_16504);
  or g48682 (n_19097, n_16417, wc1080);
  not gc1080 (wc1080, n_19093);
  or g48683 (n_18243, n_18242, wc1081);
  not gc1081 (wc1081, n_16356);
  or g48684 (n_17020, n_18577, wc1082);
  not gc1082 (wc1082, data_stack_pointer[0]);
  or g48685 (n_17008, n_18574, wc1083);
  not gc1083 (wc1083, data_stack_pointer[0]);
  or g48686 (n_18456, n_18455, wc1084);
  not gc1084 (wc1084, data_stack_pointer[0]);
  or g48687 (n_17733, wc1085, n_17944);
  not gc1085 (wc1085, n_17073);
  or g48688 (n_19462, n_19461, wc1086);
  not gc1086 (wc1086, n_17265);
  or g48689 (n_16380, wc1087, n_18301);
  not gc1087 (wc1087, n_16360);
  or g48690 (n_18347, n_18346, wc1088);
  not gc1088 (wc1088, n_16162);
  or g48691 (n_16405, wc1089, n_18313);
  not gc1089 (wc1089, n_16360);
  or g48692 (n_18324, n_18322, wc1090);
  not gc1090 (wc1090, n_16162);
  or g48693 (n_18200, n_18199, wc1091);
  not gc1091 (wc1091, n_16281);
  or g48694 (n_18179, n_18178, wc1092);
  not gc1092 (wc1092, n_16436);
  or g48695 (n_18521, wc1093, n_18518);
  not gc1093 (wc1093, n_18517);
  or g48696 (n_18223, n_18222, wc1094);
  not gc1094 (wc1094, n_16157);
  or g48697 (n_18082, n_18081, wc1095);
  not gc1095 (wc1095, n_16778);
  or g48698 (n_18146, n_18145, wc1096);
  not gc1096 (wc1096, n_16212);
  or g48699 (n_18125, n_18124, wc1097);
  not gc1097 (wc1097, n_16603);
  or g48700 (n_18064, n_18063, wc1098);
  not gc1098 (wc1098, n_16505);
  or g48701 (n_18244, n_18243, wc1099);
  not gc1099 (wc1099, n_16357);
  or g48702 (n_16986, wc1100, n_18568);
  not gc1100 (wc1100, n_16133);
  or g48703 (n_24647, wc1101, sh_reg_in[0]);
  not gc1101 (wc1101, n_16944);
  or g48704 (n_24648, n_16944, wc1102);
  not gc1102 (wc1102, sh_reg_in[0]);
  or g48705 (n_23022, n_23021, wc1103);
  not gc1103 (wc1103, data_stack_pointer[3]);
  or g48706 (n_17654, n_18913, wc1104);
  not gc1104 (wc1104, n_16160);
  or g48707 (n_23032, wc1105, n_16557);
  not gc1105 (wc1105, n_16521);
  or g48708 (n_23034, n_16522, wc1106);
  not gc1106 (wc1106, n_16557);
  or g48709 (n_16144, wc1107, n_16108);
  not gc1107 (wc1107, n_16143);
  or g48710 (n_24574, wc1108, n_16277);
  not gc1108 (wc1108, n_16267);
  or g48711 (n_24575, n_16267, wc1109);
  not gc1109 (wc1109, n_16277);
  or g48712 (n_18201, n_18200, wc1110);
  not gc1110 (wc1110, n_16268);
  or g48713 (n_24576, wc1111, n_16442);
  not gc1111 (wc1111, n_16432);
  or g48714 (n_24577, n_16432, wc1112);
  not gc1112 (wc1112, n_16442);
  or g48715 (n_18180, n_18179, wc1113);
  not gc1113 (wc1113, n_16446);
  or g48716 (n_18224, n_18223, wc1114);
  not gc1114 (wc1114, n_16159);
  or g48717 (n_24580, wc1115, n_16782);
  not gc1115 (wc1115, n_16776);
  or g48718 (n_24581, n_16776, wc1116);
  not gc1116 (wc1116, n_16782);
  or g48719 (n_18083, n_18082, wc1117);
  not gc1117 (wc1117, n_17467);
  or g48720 (n_18147, n_18146, wc1118);
  not gc1118 (wc1118, n_16200);
  or g48721 (n_24570, wc1119, n_16599);
  not gc1119 (wc1119, n_16589);
  or g48722 (n_24571, n_16589, wc1120);
  not gc1120 (wc1120, n_16599);
  or g48723 (n_18126, n_18125, wc1121);
  not gc1121 (wc1121, n_16593);
  or g48724 (n_16500, n_18034, wc1122);
  not gc1122 (wc1122, \data_stack_mem[0] [5]);
  or g48725 (n_16507, n_18064, wc1123);
  not gc1123 (wc1123, n_16506);
  or g48726 (n_24578, wc1124, n_16364);
  not gc1124 (wc1124, n_16363);
  or g48727 (n_24579, n_16363, wc1125);
  not gc1125 (wc1125, n_16364);
  or g48728 (n_18245, n_18244, wc1126);
  not gc1126 (wc1126, n_16367);
  or g48729 (n_16951, wc1127, n_18559);
  not gc1127 (wc1127, n_16133);
  or g48730 (n_17032, n_16986, wc1128);
  not gc1128 (wc1128, n_19147);
  or g48731 (n_16987, n_16986, wc1129);
  not gc1129 (wc1129, n_19150);
  or g48732 (n_18609, wc1130, n_16119);
  not gc1130 (wc1130, n_16108);
  or g48733 (n_18615, wc1131, n_16122);
  not gc1131 (wc1131, n_16108);
  or g48734 (n_18621, wc1132, n_16125);
  not gc1132 (wc1132, n_16108);
  or g48735 (n_18627, wc1133, n_16128);
  not gc1133 (wc1133, n_16108);
  or g48736 (n_18633, wc1134, n_16131);
  not gc1134 (wc1134, n_16108);
  or g48737 (n_18591, wc1135, n_16110);
  not gc1135 (wc1135, n_16108);
  or g48738 (n_18597, wc1136, n_16113);
  not gc1136 (wc1136, n_16108);
  or g48739 (n_16484, wc1137, n_18349);
  not gc1137 (wc1137, n_16439);
  or g48740 (n_18540, n_18537, wc1138);
  not gc1138 (wc1138, n_16162);
  or g48741 (n_16460, wc1139, n_18325);
  not gc1139 (wc1139, n_16439);
  or g48742 (n_23033, n_23032, wc1140);
  not gc1140 (wc1140, n_16162);
  or g48743 (n_19041, wc1141, n_19040);
  not gc1141 (wc1141, n_16302);
  or g48744 (n_18202, n_18201, wc1142);
  not gc1142 (wc1142, n_16279);
  or g48745 (n_19011, wc1143, n_19010);
  not gc1143 (wc1143, n_16467);
  or g48746 (n_18181, n_18180, wc1144);
  not gc1144 (wc1144, n_16444);
  or g48747 (n_18225, n_18224, wc1145);
  not gc1145 (wc1145, n_16161);
  or g48748 (n_19071, wc1146, n_19070);
  not gc1146 (wc1146, n_16690);
  or g48749 (n_18084, n_18083, wc1147);
  not gc1147 (wc1147, n_16667);
  or g48750 (n_18982, wc1148, n_18981);
  not gc1148 (wc1148, n_16235);
  or g48751 (n_18148, n_18147, wc1149);
  not gc1149 (wc1149, n_16210);
  or g48752 (n_18948, wc1150, n_18947);
  not gc1150 (wc1150, n_16624);
  or g48753 (n_18127, n_18126, wc1151);
  not gc1151 (wc1151, n_16601);
  or g48754 (n_19101, wc1152, n_19100);
  not gc1152 (wc1152, n_17260);
  or g48755 (n_18246, n_18245, wc1153);
  not gc1153 (wc1153, n_16353);
  or g48756 (n_16952, n_16951, wc1154);
  not gc1154 (wc1154, n_19132);
  or g48757 (n_19925, wc1155, n_19921);
  not gc1155 (wc1155, n_19920);
  or g48758 (n_20501, wc1156, n_20497);
  not gc1156 (wc1156, n_20496);
  or g48759 (n_19685, wc1157, n_19681);
  not gc1157 (wc1157, n_19680);
  or g48760 (n_24636, wc1158, n_16945);
  not gc1158 (wc1158, n_16940);
  or g48761 (n_24637, n_16940, wc1159);
  not gc1159 (wc1159, n_16945);
  or g48762 (n_20549, wc1160, n_20545);
  not gc1160 (wc1160, n_20544);
  or g48763 (n_19781, wc1161, n_19777);
  not gc1161 (wc1161, n_19776);
  or g48764 (n_16963, n_16951, wc1162);
  not gc1162 (wc1162, n_19135);
  or g48765 (n_20117, wc1163, n_20113);
  not gc1163 (wc1163, n_20112);
  or g48766 (n_20645, wc1164, n_20641);
  not gc1164 (wc1164, n_20640);
  or g48767 (n_20405, wc1165, n_20401);
  not gc1165 (wc1165, n_20400);
  or g48768 (n_19877, wc1166, n_19873);
  not gc1166 (wc1166, n_19872);
  or g48769 (n_20597, wc1167, n_20593);
  not gc1167 (wc1167, n_20592);
  or g48770 (n_20453, wc1168, n_20449);
  not gc1168 (wc1168, n_20448);
  or g48771 (n_20021, wc1169, n_20017);
  not gc1169 (wc1169, n_20016);
  or g48772 (n_20069, wc1170, n_20065);
  not gc1170 (wc1170, n_20064);
  or g48773 (n_20693, wc1171, n_20689);
  not gc1171 (wc1171, n_20688);
  or g48774 (n_19733, wc1172, n_19729);
  not gc1172 (wc1172, n_19728);
  or g48775 (n_20309, wc1173, n_20305);
  not gc1173 (wc1173, n_20304);
  or g48776 (n_19829, wc1174, n_19825);
  not gc1174 (wc1174, n_19824);
  or g48777 (n_20261, wc1175, n_20257);
  not gc1175 (wc1175, n_20256);
  or g48778 (n_20357, wc1176, n_20353);
  not gc1176 (wc1176, n_20352);
  or g48779 (n_19973, wc1177, n_19969);
  not gc1177 (wc1177, n_19968);
  or g48780 (n_20213, wc1178, n_20209);
  not gc1178 (wc1178, n_20208);
  or g48781 (n_20165, wc1179, n_20161);
  not gc1179 (wc1179, n_20160);
  or g48782 (n_16223, n_19591, wc1180);
  not gc1180 (wc1180, n_16158);
  or g48783 (n_16524, wc1181, n_18541);
  not gc1181 (wc1181, n_18540);
  or g48784 (n_19128, n_16595, wc1182);
  not gc1182 (wc1182, n_16643);
  or g48785 (n_16248, n_19597, wc1183);
  not gc1183 (wc1183, n_16158);
  or g48786 (n_19114, n_16594, wc1184);
  not gc1184 (wc1184, n_16617);
  or g48787 (n_24553, wc1185, n_16279);
  not gc1185 (wc1185, n_16278);
  or g48788 (n_24554, n_16278, wc1186);
  not gc1186 (wc1186, n_16279);
  or g48789 (n_24555, wc1187, n_16444);
  not gc1187 (wc1187, n_16443);
  or g48790 (n_24556, n_16443, wc1188);
  not gc1188 (wc1188, n_16444);
  or g48791 (n_18226, n_18225, wc1189);
  not gc1189 (wc1189, n_16149);
  or g48792 (n_24551, wc1190, n_16783);
  not gc1190 (wc1190, n_16773);
  or g48793 (n_24552, n_16773, wc1191);
  not gc1191 (wc1191, n_16783);
  or g48794 (n_18085, n_18084, wc1192);
  not gc1192 (wc1192, n_16676);
  or g48795 (n_24564, wc1193, n_16208);
  not gc1193 (wc1193, n_16198);
  or g48796 (n_24565, n_16198, wc1194);
  not gc1194 (wc1194, n_16208);
  or g48797 (n_24557, wc1195, n_16601);
  not gc1195 (wc1195, n_16600);
  or g48798 (n_24558, n_16600, wc1196);
  not gc1196 (wc1196, n_16601);
  or g48799 (n_18247, n_18246, wc1197);
  not gc1197 (wc1197, n_16364);
  or g48800 (n_18729, n_16131, wc1198);
  not gc1198 (wc1198, n_16907);
  or g48801 (n_18723, n_16128, wc1199);
  not gc1199 (wc1199, n_16907);
  or g48802 (n_18717, n_16125, wc1200);
  not gc1200 (wc1200, n_16907);
  or g48803 (n_18711, n_16122, wc1201);
  not gc1201 (wc1201, n_16907);
  or g48804 (n_18705, n_16119, wc1202);
  not gc1202 (wc1202, n_16907);
  or g48805 (n_18699, n_16116, wc1203);
  not gc1203 (wc1203, n_16907);
  or g48806 (n_18693, n_16113, wc1204);
  not gc1204 (wc1204, n_16907);
  or g48807 (n_18687, n_16110, wc1205);
  not gc1205 (wc1205, n_16907);
  or g48808 (n_16292, n_20719, wc1206);
  not gc1206 (wc1206, n_16160);
  or g48809 (n_19127, n_19126, wc1207);
  not gc1207 (wc1207, n_16162);
  or g48810 (n_16318, n_20725, wc1208);
  not gc1208 (wc1208, n_16160);
  or g48811 (n_16558, wc1209, n_23035);
  not gc1209 (wc1209, n_18539);
  or g48812 (n_19116, n_19114, wc1210);
  not gc1210 (wc1210, n_16162);
  or g48813 (n_18487, n_16507, wc1211);
  not gc1211 (wc1211, n_17751);
  or g48814 (n_19203, wc1212, n_16950);
  not gc1212 (wc1212, n_16946);
  or g48815 (n_19365, wc1213, n_16997);
  not gc1213 (wc1213, n_16946);
  or g48816 (n_19257, wc1214, n_16962);
  not gc1214 (wc1214, n_16946);
  or g48817 (n_19389, wc1215, n_17031);
  not gc1215 (wc1215, n_16946);
  or g48818 (n_19287, wc1216, n_16985);
  not gc1216 (wc1216, n_16946);
  or g48819 (n_18891, wc1217, n_16973);
  not gc1217 (wc1217, n_16946);
  or g48820 (n_18837, wc1218, n_17042);
  not gc1218 (wc1218, n_16946);
  or g48821 (n_18831, wc1219, n_16927);
  not gc1219 (wc1219, n_16946);
  or g48822 (n_19437, n_16681, wc1220);
  not gc1220 (wc1220, n_16683);
  or g48823 (n_19447, n_16680, wc1221);
  not gc1221 (wc1221, n_16731);
  or g48824 (n_23014, n_17467, wc1222);
  not gc1222 (wc1222, n_16731);
  or g48825 (n_24541, wc1223, n_16281);
  not gc1223 (wc1223, n_16280);
  or g48826 (n_24542, n_16280, wc1224);
  not gc1224 (wc1224, n_16281);
  or g48827 (n_24537, wc1225, n_16446);
  not gc1225 (wc1225, n_16445);
  or g48828 (n_24538, n_16445, wc1226);
  not gc1226 (wc1226, n_16446);
  or g48829 (n_24545, wc1227, n_16210);
  not gc1227 (wc1227, n_16209);
  or g48830 (n_24546, n_16209, wc1228);
  not gc1228 (wc1228, n_16210);
  or g48831 (n_24535, wc1229, n_16603);
  not gc1229 (wc1229, n_16602);
  or g48832 (n_24536, n_16602, wc1230);
  not gc1230 (wc1230, n_16603);
  or g48833 (n_16644, wc1231, n_19129);
  not gc1231 (wc1231, n_16596);
  or g48834 (n_19436, n_19435, wc1232);
  not gc1232 (wc1232, n_16162);
  or g48835 (n_16618, wc1233, n_19117);
  not gc1233 (wc1233, n_16596);
  or g48836 (n_19449, n_19447, wc1234);
  not gc1234 (wc1234, n_16162);
  or g48837 (n_16378, n_20809, wc1235);
  not gc1235 (wc1235, n_16160);
  or g48838 (n_20925, n_16321, wc1236);
  not gc1236 (wc1236, n_17642);
  or g48839 (n_20926, wc1237, n_17642);
  not gc1237 (wc1237, n_16321);
  or g48840 (n_16403, n_20815, wc1238);
  not gc1238 (wc1238, n_16160);
  or g48841 (n_24529, wc1239, n_16212);
  not gc1239 (wc1239, n_16211);
  or g48842 (n_24530, n_16211, wc1240);
  not gc1240 (wc1240, n_16212);
  or g48843 (n_24531, wc1241, n_16368);
  not gc1241 (wc1241, n_16354);
  or g48844 (n_24532, n_16354, wc1242);
  not gc1242 (wc1242, n_16368);
  or g48845 (n_20862, n_16295, wc1243);
  not gc1243 (wc1243, n_17653);
  or g48846 (n_20863, wc1244, n_17653);
  not gc1244 (wc1244, n_16295);
  or g48847 (n_16684, wc1245, n_19438);
  not gc1245 (wc1245, n_16682);
  or g48848 (n_16732, wc1246, n_19450);
  not gc1246 (wc1246, n_16682);
  or g48849 (n_16217, n_20797, wc1247);
  not gc1247 (wc1247, n_16152);
  or g48850 (n_21017, n_21015, wc1248);
  not gc1248 (wc1248, n_16160);
  or g48851 (n_16242, n_20803, wc1249);
  not gc1249 (wc1249, n_16152);
  or g48852 (n_17669, n_20896, wc1250);
  not gc1250 (wc1250, n_16160);
  or g48853 (n_17672, n_20974, wc1251);
  not gc1251 (wc1251, n_16160);
  or g48854 (n_21078, n_16381, wc1252);
  not gc1252 (wc1252, n_17657);
  or g48855 (n_21079, wc1253, n_17657);
  not gc1253 (wc1253, n_16381);
  or g48856 (n_21072, n_16406, wc1254);
  not gc1254 (wc1254, n_17650);
  or g48857 (n_21073, wc1255, n_17650);
  not gc1255 (wc1255, n_16406);
  or g48858 (n_17674, n_20830, wc1256);
  not gc1256 (wc1256, n_16148);
  or g48859 (n_16520, n_21043, wc1257);
  not gc1257 (wc1257, n_16160);
  or g48860 (n_20998, n_16171, wc1258);
  not gc1258 (wc1258, n_17725);
  or g48861 (n_16556, n_21184, wc1259);
  not gc1259 (wc1259, n_16160);
  or g48862 (n_16286, n_21031, wc1260);
  not gc1260 (wc1260, n_16152);
  or g48863 (n_16481, n_21178, wc1261);
  not gc1261 (wc1261, n_16158);
  or g48864 (n_16457, n_21172, wc1262);
  not gc1262 (wc1262, n_16158);
  or g48865 (n_16312, n_21037, wc1263);
  not gc1263 (wc1263, n_16152);
  or g48866 (n_17726, wc1264, n_21001);
  not gc1264 (wc1264, n_21000);
  or g48867 (n_16256, wc1265, n_21103);
  not gc1265 (wc1265, n_21102);
  or g48868 (n_21112, wc1266, n_16185);
  not gc1266 (wc1266, n_17726);
  or g48869 (n_16518, n_21304, wc1267);
  not gc1267 (wc1267, n_16158);
  or g48870 (n_16554, n_21298, wc1268);
  not gc1268 (wc1268, n_16158);
  or g48871 (n_17665, n_21193, wc1269);
  not gc1269 (wc1269, n_16148);
  or g48872 (n_16373, n_21286, wc1270);
  not gc1270 (wc1270, n_16152);
  or g48873 (n_16397, n_21292, wc1271);
  not gc1271 (wc1271, n_16152);
  or g48874 (n_16641, n_21490, wc1272);
  not gc1272 (wc1272, n_16158);
  or g48875 (n_16614, n_21484, wc1273);
  not gc1273 (wc1273, n_16158);
  or g48876 (n_16328, wc1274, n_21355);
  not gc1274 (wc1274, n_21354);
  or g48877 (n_21436, n_17260, wc1275);
  not gc1275 (wc1275, n_16412);
  or g48878 (n_21337, n_16306, wc1276);
  not gc1276 (wc1276, n_16330);
  or g48879 (n_16746, n_17448, wc1277);
  not gc1277 (wc1277, n_21661);
  or g48880 (n_16477, n_21556, wc1278);
  not gc1278 (wc1278, n_16152);
  or g48881 (n_16451, n_21550, wc1279);
  not gc1279 (wc1279, n_16152);
  or g48882 (n_21862, n_16800, wc1280);
  not gc1280 (wc1280, n_16701);
  or g48883 (n_21517, wc1281, n_21516);
  not gc1281 (wc1281, n_21515);
  or g48884 (n_16262, n_16144, wc1282);
  not gc1282 (wc1282, n_21376);
  or g48885 (n_21817, n_16734, wc1283);
  not gc1283 (wc1283, n_17336);
  or g48886 (n_17644, n_21565, wc1284);
  not gc1284 (wc1284, n_16148);
  or g48887 (n_16697, n_17335, wc1285);
  not gc1285 (wc1285, n_21841);
  or g48888 (n_16548, n_21778, wc1286);
  not gc1286 (wc1286, n_16152);
  or g48889 (n_21595, wc1287, n_21594);
  not gc1287 (wc1287, n_21593);
  or g48890 (n_21658, n_16391, wc1288);
  not gc1288 (wc1288, n_16415);
  or g48891 (n_17382, n_21733, wc1289);
  not gc1289 (wc1289, n_16152);
  or g48892 (n_16817, n_16745, wc1290);
  not gc1290 (wc1290, n_16750);
  or g48893 (n_17287, n_16817, wc1291);
  not gc1291 (wc1291, n_16820);
  or g48894 (n_21748, wc1292, n_21747);
  not gc1292 (wc1292, n_21746);
  or g48895 (n_21801, n_16414, wc1293);
  not gc1293 (wc1293, n_17698);
  or g48896 (n_21967, n_16735, wc1294);
  not gc1294 (wc1294, n_17318);
  or g48897 (n_16469, wc1295, n_21832);
  not gc1295 (wc1295, n_21831);
  or g48898 (n_16511, n_21847, wc1296);
  not gc1296 (wc1296, n_16148);
  or g48899 (n_16635, n_21931, wc1297);
  not gc1297 (wc1297, n_16152);
  or g48900 (n_16608, n_21925, wc1298);
  not gc1298 (wc1298, n_16152);
  or g48901 (n_16335, n_16144, wc1299);
  not gc1299 (wc1299, n_21673);
  or g48902 (n_21961, n_16471, wc1300);
  not gc1300 (wc1300, n_16492);
  or g48903 (n_21805, wc1301, n_21804);
  not gc1301 (wc1301, n_21803);
  or g48904 (n_16816, n_16744, wc1302);
  not gc1302 (wc1302, n_16751);
  or g48905 (n_16546, n_21937, wc1303);
  not gc1303 (wc1303, n_16148);
  or g48906 (n_21988, n_16624, wc1304);
  not gc1304 (wc1304, n_16625);
  or g48907 (n_17371, n_16816, wc1305);
  not gc1305 (wc1305, n_16821);
  or g48908 (n_22002, n_16493, wc1306);
  not gc1306 (wc1306, n_17696);
  or g48909 (n_22051, n_16736, wc1307);
  not gc1307 (wc1307, n_17454);
  or g48910 (n_17651, n_21952, wc1308);
  not gc1308 (wc1308, n_16148);
  or g48911 (n_16708, n_17453, wc1309);
  not gc1309 (wc1309, n_22054);
  or g48912 (n_22098, n_16623, wc1310);
  not gc1310 (wc1310, n_17638);
  or g48913 (n_22099, wc1311, n_17638);
  not gc1311 (wc1311, n_16623);
  or g48914 (n_22006, wc1312, n_22005);
  not gc1312 (wc1312, n_22004);
  or g48915 (n_22041, n_16472, wc1313);
  not gc1313 (wc1313, n_17693);
  or g48916 (n_16420, n_16144, wc1314);
  not gc1314 (wc1314, n_21871);
  or g48917 (n_16815, n_16743, wc1315);
  not gc1315 (wc1315, n_16752);
  or g48918 (n_22072, n_16690, wc1316);
  not gc1316 (wc1316, n_16738);
  or g48919 (n_17354, n_16815, wc1317);
  not gc1317 (wc1317, n_16822);
  or g48920 (n_22045, wc1318, n_22044);
  not gc1318 (wc1318, n_22043);
  or g48921 (n_22085, n_16531, wc1319);
  not gc1319 (wc1319, n_16533);
  or g48922 (n_22086, wc1320, n_16533);
  not gc1320 (wc1320, n_16531);
  or g48923 (n_22219, n_16737, wc1321);
  not gc1321 (wc1321, n_17462);
  or g48924 (n_22248, n_16737, wc1322);
  not gc1322 (wc1322, n_17647);
  or g48925 (n_22249, wc1323, n_17647);
  not gc1323 (wc1323, n_16737);
  or g48926 (n_24351, wc1324, n_16806);
  not gc1324 (wc1324, n_16801);
  or g48927 (n_24352, n_16801, wc1325);
  not gc1325 (wc1325, n_16806);
  or g48928 (n_22278, n_16689, wc1326);
  not gc1326 (wc1326, n_17658);
  or g48929 (n_22279, wc1327, n_17658);
  not gc1327 (wc1327, n_16689);
  or g48930 (n_16695, n_16692, wc1328);
  not gc1328 (wc1328, n_22252);
  or g48931 (n_22184, wc1329, n_16567);
  not gc1329 (wc1329, n_16565);
  or g48932 (n_22185, n_16565, wc1330);
  not gc1330 (wc1330, n_16567);
  or g48933 (n_16814, n_16742, wc1331);
  not gc1331 (wc1331, n_16753);
  or g48934 (n_24339, wc1332, n_16804);
  not gc1332 (wc1332, n_16807);
  or g48935 (n_24340, n_16807, wc1333);
  not gc1333 (wc1333, n_16804);
  or g48936 (n_22204, n_16628, wc1334);
  not gc1334 (wc1334, n_16629);
  or g48937 (n_16498, n_16144, wc1335);
  not gc1335 (wc1335, n_22129);
  or g48938 (n_16829, wc1336, n_16828);
  not gc1336 (wc1336, n_17440);
  or g48939 (n_24329, wc1337, n_16810);
  not gc1337 (wc1337, n_16808);
  or g48940 (n_24330, n_16808, wc1338);
  not gc1338 (wc1338, n_16810);
  or g48941 (n_16825, wc1339, n_16741);
  not gc1339 (wc1339, n_16754);
  or g48942 (n_22418, n_16801, wc1340);
  not gc1340 (wc1340, n_16694);
  or g48943 (n_22284, wc1341, n_16569);
  not gc1341 (wc1341, n_17690);
  or g48944 (n_22419, n_22418, wc1342);
  not gc1342 (wc1342, n_16696);
  or g48945 (n_24323, wc1343, n_16812);
  not gc1343 (wc1343, n_17284);
  or g48946 (n_24324, n_17284, wc1344);
  not gc1344 (wc1344, n_16812);
  or g48947 (n_22420, n_22419, wc1345);
  not gc1345 (wc1345, n_16708);
  or g48948 (n_22446, wc1346, n_16771);
  not gc1346 (wc1346, n_16757);
  or g48949 (n_16570, n_16144, wc1347);
  not gc1347 (wc1347, n_22285);
  or g48950 (n_16719, n_16718, wc1348);
  not gc1348 (wc1348, n_22423);
  or g48951 (n_16850, n_22420, wc1349);
  not gc1349 (wc1349, n_16695);
  or g48952 (n_22428, n_16850, wc1350);
  not gc1350 (wc1350, n_16719);
  or g48953 (n_22463, n_16719, wc1351);
  not gc1351 (wc1351, n_16714);
  or g48954 (n_22464, wc1352, n_16714);
  not gc1352 (wc1352, n_16719);
  or g48955 (n_16657, n_16144, wc1353);
  not gc1353 (wc1353, n_22351);
  or g48956 (n_22429, wc1354, n_16144);
  not gc1354 (wc1354, n_22428);
  or g48957 (n_16760, n_17439, wc1355);
  not gc1355 (wc1355, n_16755);
  or g48958 (n_22638, n_16755, wc1356);
  not gc1356 (wc1356, n_17439);
  or g48959 (n_16833, wc1357, n_16832);
  not gc1357 (wc1357, n_16830);
  or g48960 (n_22773, n_16830, wc1358);
  not gc1358 (wc1358, n_16832);
  or g48961 (n_16791, n_16144, wc1359);
  not gc1359 (wc1359, n_22480);
  or g48962 (n_16762, n_16144, wc1360);
  not gc1360 (wc1360, n_22672);
  or g48963 (n_16848, n_16144, wc1361);
  not gc1361 (wc1361, n_22669);
  or g48964 (n_16852, n_16144, wc1362);
  not gc1362 (wc1362, n_22834);
  or g48965 (n_16838, n_16144, wc1363);
  not gc1363 (wc1363, n_22837);
  or g48966 (n_22785, n_16113, wc1364);
  not gc1364 (wc1364, n_16874);
  or g48967 (n_22791, n_16116, wc1365);
  not gc1365 (wc1365, n_16874);
  or g48968 (n_22779, n_16110, wc1366);
  not gc1366 (wc1366, n_16874);
  or g48969 (n_22797, n_16119, wc1367);
  not gc1367 (wc1367, n_16874);
  or g48970 (n_22803, n_16122, wc1368);
  not gc1368 (wc1368, n_16874);
  or g48971 (n_22809, n_16125, wc1369);
  not gc1369 (wc1369, n_16874);
  or g48972 (n_22821, n_16131, wc1370);
  not gc1370 (wc1370, n_16874);
  or g48973 (n_22815, n_16128, wc1371);
  not gc1371 (wc1371, n_16874);
  or g48974 (n_22938, n_16110, wc1372);
  not gc1372 (wc1372, n_16889);
  or g48975 (n_22944, n_16113, wc1373);
  not gc1373 (wc1373, n_16889);
  or g48976 (n_22950, n_16116, wc1374);
  not gc1374 (wc1374, n_16889);
  or g48977 (n_22980, n_16131, wc1375);
  not gc1375 (wc1375, n_16889);
  or g48978 (n_22962, n_16122, wc1376);
  not gc1376 (wc1376, n_16889);
  or g48979 (n_22968, n_16125, wc1377);
  not gc1377 (wc1377, n_16889);
  or g48980 (n_22974, n_16128, wc1378);
  not gc1378 (wc1378, n_16889);
  or g48981 (n_22956, n_16119, wc1379);
  not gc1379 (wc1379, n_16889);
  CDN_flop \out_fifo_read_pointer_reg[0] (.clk (clk), .d (n_24622),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[0]));
  CDN_flop \out_fifo_read_pointer_reg[1] (.clk (clk), .d (n_24596),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[1]));
  CDN_flop \out_fifo_read_pointer_reg[2] (.clk (clk), .d (n_24561),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_read_pointer[2]));
  CDN_flop \out_fifo_reg[0][0][0] (.clk (clk), .d (n_16879), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [0]));
  CDN_flop \out_fifo_reg[0][0][1] (.clk (clk), .d (n_16191), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [1]));
  CDN_flop \out_fifo_reg[0][0][2] (.clk (clk), .d (n_16343), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [2]));
  CDN_flop \out_fifo_reg[0][0][3] (.clk (clk), .d (n_16344), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [3]));
  CDN_flop \out_fifo_reg[0][0][4] (.clk (clk), .d (n_16425), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [4]));
  CDN_flop \out_fifo_reg[0][0][5] (.clk (clk), .d (n_16578), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [5]));
  CDN_flop \out_fifo_reg[0][0][6] (.clk (clk), .d (n_16579), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [6]));
  CDN_flop \out_fifo_reg[0][0][7] (.clk (clk), .d (n_16662), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [7]));
  CDN_flop \out_fifo_reg[0][0][8] (.clk (clk), .d (n_16796), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][0] [8]));
  CDN_flop \out_fifo_reg[0][1][0] (.clk (clk), .d (n_16894), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [0]));
  CDN_flop \out_fifo_reg[0][1][1] (.clk (clk), .d (n_16767), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [1]));
  CDN_flop \out_fifo_reg[0][1][2] (.clk (clk), .d (n_16860), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [2]));
  CDN_flop \out_fifo_reg[0][1][3] (.clk (clk), .d (n_16843), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [3]));
  CDN_flop \out_fifo_reg[0][1][4] (.clk (clk), .d (n_16861), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [4]));
  CDN_flop \out_fifo_reg[0][1][5] (.clk (clk), .d (n_17101), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [5]));
  CDN_flop \out_fifo_reg[0][1][6] (.clk (clk), .d (n_17098), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [6]));
  CDN_flop \out_fifo_reg[0][1][7] (.clk (clk), .d (n_17099), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [7]));
  CDN_flop \out_fifo_reg[0][1][8] (.clk (clk), .d (n_17100), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][1] [8]));
  CDN_flop \out_fifo_reg[0][2][0] (.clk (clk), .d (n_16912), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [0]));
  CDN_flop \out_fifo_reg[0][2][1] (.clk (clk), .d (n_16920), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [1]));
  CDN_flop \out_fifo_reg[0][2][6] (.clk (clk), .d (n_16123), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [6]));
  CDN_flop \out_fifo_reg[0][2][8] (.clk (clk), .d (n_16903), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[0][2] [8]));
  CDN_flop \out_fifo_reg[0][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16095), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (\out_fifo[0][2] [9]));
  CDN_flop \out_fifo_reg[1][0][0] (.clk (clk), .d (n_16882), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [0]));
  CDN_flop \out_fifo_reg[1][0][1] (.clk (clk), .d (n_16194), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [1]));
  CDN_flop \out_fifo_reg[1][0][2] (.clk (clk), .d (n_16349), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [2]));
  CDN_flop \out_fifo_reg[1][0][3] (.clk (clk), .d (n_16350), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [3]));
  CDN_flop \out_fifo_reg[1][0][4] (.clk (clk), .d (n_16428), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [4]));
  CDN_flop \out_fifo_reg[1][0][5] (.clk (clk), .d (n_16584), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [5]));
  CDN_flop \out_fifo_reg[1][0][6] (.clk (clk), .d (n_16585), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [6]));
  CDN_flop \out_fifo_reg[1][0][7] (.clk (clk), .d (n_16665), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [7]));
  CDN_flop \out_fifo_reg[1][0][8] (.clk (clk), .d (n_16799), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][0] [8]));
  CDN_flop \out_fifo_reg[1][1][0] (.clk (clk), .d (n_16897), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [0]));
  CDN_flop \out_fifo_reg[1][1][1] (.clk (clk), .d (n_16770), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [1]));
  CDN_flop \out_fifo_reg[1][1][2] (.clk (clk), .d (n_16866), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [2]));
  CDN_flop \out_fifo_reg[1][1][3] (.clk (clk), .d (n_16846), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [3]));
  CDN_flop \out_fifo_reg[1][1][4] (.clk (clk), .d (n_16867), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [4]));
  CDN_flop \out_fifo_reg[1][1][5] (.clk (clk), .d (n_17088), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [5]));
  CDN_flop \out_fifo_reg[1][1][6] (.clk (clk), .d (n_17089), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [6]));
  CDN_flop \out_fifo_reg[1][1][7] (.clk (clk), .d (n_17090), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [7]));
  CDN_flop \out_fifo_reg[1][1][8] (.clk (clk), .d (n_17091), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][1] [8]));
  CDN_flop \out_fifo_reg[1][2][0] (.clk (clk), .d (n_16915), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [0]));
  CDN_flop \out_fifo_reg[1][2][1] (.clk (clk), .d (n_16923), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [1]));
  CDN_flop \out_fifo_reg[1][2][6] (.clk (clk), .d (n_16132), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [6]));
  CDN_flop \out_fifo_reg[1][2][8] (.clk (clk), .d (n_16906), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[1][2] [8]));
  CDN_flop \out_fifo_reg[1][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16093), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (\out_fifo[1][2] [9]));
  CDN_flop \out_fifo_reg[2][0][0] (.clk (clk), .d (n_16880), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [0]));
  CDN_flop \out_fifo_reg[2][0][1] (.clk (clk), .d (n_16192), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [1]));
  CDN_flop \out_fifo_reg[2][0][2] (.clk (clk), .d (n_16345), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [2]));
  CDN_flop \out_fifo_reg[2][0][3] (.clk (clk), .d (n_16346), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [3]));
  CDN_flop \out_fifo_reg[2][0][4] (.clk (clk), .d (n_16426), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [4]));
  CDN_flop \out_fifo_reg[2][0][5] (.clk (clk), .d (n_16580), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [5]));
  CDN_flop \out_fifo_reg[2][0][6] (.clk (clk), .d (n_16581), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [6]));
  CDN_flop \out_fifo_reg[2][0][7] (.clk (clk), .d (n_16663), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [7]));
  CDN_flop \out_fifo_reg[2][0][8] (.clk (clk), .d (n_16797), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][0] [8]));
  CDN_flop \out_fifo_reg[2][1][0] (.clk (clk), .d (n_16895), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [0]));
  CDN_flop \out_fifo_reg[2][1][1] (.clk (clk), .d (n_16768), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [1]));
  CDN_flop \out_fifo_reg[2][1][2] (.clk (clk), .d (n_16862), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [2]));
  CDN_flop \out_fifo_reg[2][1][3] (.clk (clk), .d (n_16844), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [3]));
  CDN_flop \out_fifo_reg[2][1][4] (.clk (clk), .d (n_16863), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [4]));
  CDN_flop \out_fifo_reg[2][1][5] (.clk (clk), .d (n_17095), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [5]));
  CDN_flop \out_fifo_reg[2][1][6] (.clk (clk), .d (n_17093), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [6]));
  CDN_flop \out_fifo_reg[2][1][7] (.clk (clk), .d (n_17096), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [7]));
  CDN_flop \out_fifo_reg[2][1][8] (.clk (clk), .d (n_17094), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][1] [8]));
  CDN_flop \out_fifo_reg[2][2][0] (.clk (clk), .d (n_16913), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [0]));
  CDN_flop \out_fifo_reg[2][2][1] (.clk (clk), .d (n_16921), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [1]));
  CDN_flop \out_fifo_reg[2][2][6] (.clk (clk), .d (n_16126), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [6]));
  CDN_flop \out_fifo_reg[2][2][8] (.clk (clk), .d (n_16904), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[2][2] [8]));
  CDN_flop \out_fifo_reg[2][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16091), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (\out_fifo[2][2] [9]));
  CDN_flop \out_fifo_reg[3][0][0] (.clk (clk), .d (n_16877), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [0]));
  CDN_flop \out_fifo_reg[3][0][1] (.clk (clk), .d (n_16189), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [1]));
  CDN_flop \out_fifo_reg[3][0][2] (.clk (clk), .d (n_16339), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [2]));
  CDN_flop \out_fifo_reg[3][0][3] (.clk (clk), .d (n_16340), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [3]));
  CDN_flop \out_fifo_reg[3][0][4] (.clk (clk), .d (n_16423), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [4]));
  CDN_flop \out_fifo_reg[3][0][5] (.clk (clk), .d (n_16574), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [5]));
  CDN_flop \out_fifo_reg[3][0][6] (.clk (clk), .d (n_16575), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [6]));
  CDN_flop \out_fifo_reg[3][0][7] (.clk (clk), .d (n_16660), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [7]));
  CDN_flop \out_fifo_reg[3][0][8] (.clk (clk), .d (n_16794), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][0] [8]));
  CDN_flop \out_fifo_reg[3][1][0] (.clk (clk), .d (n_16892), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [0]));
  CDN_flop \out_fifo_reg[3][1][1] (.clk (clk), .d (n_16765), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [1]));
  CDN_flop \out_fifo_reg[3][1][2] (.clk (clk), .d (n_16856), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [2]));
  CDN_flop \out_fifo_reg[3][1][3] (.clk (clk), .d (n_16841), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [3]));
  CDN_flop \out_fifo_reg[3][1][4] (.clk (clk), .d (n_16857), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [4]));
  CDN_flop \out_fifo_reg[3][1][5] (.clk (clk), .d (n_17105), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [5]));
  CDN_flop \out_fifo_reg[3][1][6] (.clk (clk), .d (n_17104), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [6]));
  CDN_flop \out_fifo_reg[3][1][7] (.clk (clk), .d (n_17103), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [7]));
  CDN_flop \out_fifo_reg[3][1][8] (.clk (clk), .d (n_17106), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][1] [8]));
  CDN_flop \out_fifo_reg[3][2][0] (.clk (clk), .d (n_16910), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [0]));
  CDN_flop \out_fifo_reg[3][2][1] (.clk (clk), .d (n_16918), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [1]));
  CDN_flop \out_fifo_reg[3][2][6] (.clk (clk), .d (n_16117), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [6]));
  CDN_flop \out_fifo_reg[3][2][8] (.clk (clk), .d (n_16901), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[3][2] [8]));
  CDN_flop \out_fifo_reg[3][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16089), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (\out_fifo[3][2] [9]));
  CDN_flop \out_fifo_reg[4][0][0] (.clk (clk), .d (n_16881), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [0]));
  CDN_flop \out_fifo_reg[4][0][1] (.clk (clk), .d (n_16193), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [1]));
  CDN_flop \out_fifo_reg[4][0][2] (.clk (clk), .d (n_16347), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [2]));
  CDN_flop \out_fifo_reg[4][0][3] (.clk (clk), .d (n_16348), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [3]));
  CDN_flop \out_fifo_reg[4][0][4] (.clk (clk), .d (n_16427), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [4]));
  CDN_flop \out_fifo_reg[4][0][5] (.clk (clk), .d (n_16582), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [5]));
  CDN_flop \out_fifo_reg[4][0][6] (.clk (clk), .d (n_16583), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [6]));
  CDN_flop \out_fifo_reg[4][0][7] (.clk (clk), .d (n_16664), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [7]));
  CDN_flop \out_fifo_reg[4][0][8] (.clk (clk), .d (n_16798), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][0] [8]));
  CDN_flop \out_fifo_reg[4][1][0] (.clk (clk), .d (n_16896), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [0]));
  CDN_flop \out_fifo_reg[4][1][1] (.clk (clk), .d (n_16769), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [1]));
  CDN_flop \out_fifo_reg[4][1][2] (.clk (clk), .d (n_16864), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [2]));
  CDN_flop \out_fifo_reg[4][1][3] (.clk (clk), .d (n_16845), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [3]));
  CDN_flop \out_fifo_reg[4][1][4] (.clk (clk), .d (n_16865), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [4]));
  CDN_flop \out_fifo_reg[4][1][5] (.clk (clk), .d (n_17121), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [5]));
  CDN_flop \out_fifo_reg[4][1][6] (.clk (clk), .d (n_17119), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [6]));
  CDN_flop \out_fifo_reg[4][1][7] (.clk (clk), .d (n_17120), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [7]));
  CDN_flop \out_fifo_reg[4][1][8] (.clk (clk), .d (n_17118), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][1] [8]));
  CDN_flop \out_fifo_reg[4][2][0] (.clk (clk), .d (n_16914), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [0]));
  CDN_flop \out_fifo_reg[4][2][1] (.clk (clk), .d (n_16922), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [1]));
  CDN_flop \out_fifo_reg[4][2][6] (.clk (clk), .d (n_16129), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [6]));
  CDN_flop \out_fifo_reg[4][2][8] (.clk (clk), .d (n_16905), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[4][2] [8]));
  CDN_flop \out_fifo_reg[4][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16087), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (\out_fifo[4][2] [9]));
  CDN_flop \out_fifo_reg[5][0][0] (.clk (clk), .d (n_16876), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [0]));
  CDN_flop \out_fifo_reg[5][0][1] (.clk (clk), .d (n_16188), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [1]));
  CDN_flop \out_fifo_reg[5][0][2] (.clk (clk), .d (n_16337), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [2]));
  CDN_flop \out_fifo_reg[5][0][3] (.clk (clk), .d (n_16338), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [3]));
  CDN_flop \out_fifo_reg[5][0][4] (.clk (clk), .d (n_16422), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [4]));
  CDN_flop \out_fifo_reg[5][0][5] (.clk (clk), .d (n_16572), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [5]));
  CDN_flop \out_fifo_reg[5][0][6] (.clk (clk), .d (n_16573), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [6]));
  CDN_flop \out_fifo_reg[5][0][7] (.clk (clk), .d (n_16659), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [7]));
  CDN_flop \out_fifo_reg[5][0][8] (.clk (clk), .d (n_16793), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][0] [8]));
  CDN_flop \out_fifo_reg[5][1][0] (.clk (clk), .d (n_16891), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [0]));
  CDN_flop \out_fifo_reg[5][1][1] (.clk (clk), .d (n_16764), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [1]));
  CDN_flop \out_fifo_reg[5][1][2] (.clk (clk), .d (n_16854), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [2]));
  CDN_flop \out_fifo_reg[5][1][3] (.clk (clk), .d (n_16840), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [3]));
  CDN_flop \out_fifo_reg[5][1][4] (.clk (clk), .d (n_16855), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [4]));
  CDN_flop \out_fifo_reg[5][1][5] (.clk (clk), .d (n_17111), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [5]));
  CDN_flop \out_fifo_reg[5][1][6] (.clk (clk), .d (n_17108), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [6]));
  CDN_flop \out_fifo_reg[5][1][7] (.clk (clk), .d (n_17109), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [7]));
  CDN_flop \out_fifo_reg[5][1][8] (.clk (clk), .d (n_17110), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][1] [8]));
  CDN_flop \out_fifo_reg[5][2][0] (.clk (clk), .d (n_16909), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [0]));
  CDN_flop \out_fifo_reg[5][2][1] (.clk (clk), .d (n_16917), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [1]));
  CDN_flop \out_fifo_reg[5][2][6] (.clk (clk), .d (n_16114), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [6]));
  CDN_flop \out_fifo_reg[5][2][8] (.clk (clk), .d (n_16900), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[5][2] [8]));
  CDN_flop \out_fifo_reg[5][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16085), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (\out_fifo[5][2] [9]));
  CDN_flop \out_fifo_reg[6][0][0] (.clk (clk), .d (n_16878), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [0]));
  CDN_flop \out_fifo_reg[6][0][1] (.clk (clk), .d (n_16190), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [1]));
  CDN_flop \out_fifo_reg[6][0][2] (.clk (clk), .d (n_16341), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [2]));
  CDN_flop \out_fifo_reg[6][0][3] (.clk (clk), .d (n_16342), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [3]));
  CDN_flop \out_fifo_reg[6][0][4] (.clk (clk), .d (n_16424), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [4]));
  CDN_flop \out_fifo_reg[6][0][5] (.clk (clk), .d (n_16576), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [5]));
  CDN_flop \out_fifo_reg[6][0][6] (.clk (clk), .d (n_16577), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [6]));
  CDN_flop \out_fifo_reg[6][0][7] (.clk (clk), .d (n_16661), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [7]));
  CDN_flop \out_fifo_reg[6][0][8] (.clk (clk), .d (n_16795), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][0] [8]));
  CDN_flop \out_fifo_reg[6][1][0] (.clk (clk), .d (n_16893), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [0]));
  CDN_flop \out_fifo_reg[6][1][1] (.clk (clk), .d (n_16766), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [1]));
  CDN_flop \out_fifo_reg[6][1][2] (.clk (clk), .d (n_16858), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [2]));
  CDN_flop \out_fifo_reg[6][1][3] (.clk (clk), .d (n_16842), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [3]));
  CDN_flop \out_fifo_reg[6][1][4] (.clk (clk), .d (n_16859), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [4]));
  CDN_flop \out_fifo_reg[6][1][5] (.clk (clk), .d (n_17114), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [5]));
  CDN_flop \out_fifo_reg[6][1][6] (.clk (clk), .d (n_17115), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [6]));
  CDN_flop \out_fifo_reg[6][1][7] (.clk (clk), .d (n_17113), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [7]));
  CDN_flop \out_fifo_reg[6][1][8] (.clk (clk), .d (n_17116), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][1] [8]));
  CDN_flop \out_fifo_reg[6][2][0] (.clk (clk), .d (n_16911), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [0]));
  CDN_flop \out_fifo_reg[6][2][1] (.clk (clk), .d (n_16919), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [1]));
  CDN_flop \out_fifo_reg[6][2][6] (.clk (clk), .d (n_16120), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [6]));
  CDN_flop \out_fifo_reg[6][2][8] (.clk (clk), .d (n_16902), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[6][2] [8]));
  CDN_flop \out_fifo_reg[6][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16082), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (\out_fifo[6][2] [9]));
  CDN_flop \out_fifo_reg[7][0][0] (.clk (clk), .d (n_16875), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [0]));
  CDN_flop \out_fifo_reg[7][0][1] (.clk (clk), .d (n_16187), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [1]));
  CDN_flop \out_fifo_reg[7][0][2] (.clk (clk), .d (n_16263), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [2]));
  CDN_flop \out_fifo_reg[7][0][3] (.clk (clk), .d (n_16336), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [3]));
  CDN_flop \out_fifo_reg[7][0][4] (.clk (clk), .d (n_16421), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [4]));
  CDN_flop \out_fifo_reg[7][0][5] (.clk (clk), .d (n_16499), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [5]));
  CDN_flop \out_fifo_reg[7][0][6] (.clk (clk), .d (n_16571), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [6]));
  CDN_flop \out_fifo_reg[7][0][7] (.clk (clk), .d (n_16658), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [7]));
  CDN_flop \out_fifo_reg[7][0][8] (.clk (clk), .d (n_16792), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][0] [8]));
  CDN_flop \out_fifo_reg[7][1][0] (.clk (clk), .d (n_16890), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [0]));
  CDN_flop \out_fifo_reg[7][1][1] (.clk (clk), .d (n_16763), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [1]));
  CDN_flop \out_fifo_reg[7][1][2] (.clk (clk), .d (n_16849), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [2]));
  CDN_flop \out_fifo_reg[7][1][3] (.clk (clk), .d (n_16839), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [3]));
  CDN_flop \out_fifo_reg[7][1][4] (.clk (clk), .d (n_16853), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [4]));
  CDN_flop \out_fifo_reg[7][1][5] (.clk (clk), .d (n_17084), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [5]));
  CDN_flop \out_fifo_reg[7][1][6] (.clk (clk), .d (n_17086), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [6]));
  CDN_flop \out_fifo_reg[7][1][7] (.clk (clk), .d (n_17085), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [7]));
  CDN_flop \out_fifo_reg[7][1][8] (.clk (clk), .d (n_17083), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][1] [8]));
  CDN_flop \out_fifo_reg[7][2][0] (.clk (clk), .d (n_16908), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [0]));
  CDN_flop \out_fifo_reg[7][2][1] (.clk (clk), .d (n_16916), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [1]));
  CDN_flop \out_fifo_reg[7][2][6] (.clk (clk), .d (n_16111), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [6]));
  CDN_flop \out_fifo_reg[7][2][8] (.clk (clk), .d (n_16899), .sena
       (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (\out_fifo[7][2] [8]));
  CDN_flop \out_fifo_reg[7][2][9] (.clk (clk), .d (1'b1), .sena
       (n_16080), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (\out_fifo[7][2] [9]));
  CDN_flop \out_fifo_write_pointer_reg[0] (.clk (clk), .d (n_24593),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[0]));
  CDN_flop \out_fifo_write_pointer_reg[1] (.clk (clk), .d (n_17056),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[1]));
  CDN_flop \out_fifo_write_pointer_reg[2] (.clk (clk), .d (n_17125),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (out_fifo_write_pointer[2]));
  CDN_flop \sh_bit_cnt_reg[0] (.clk (clk), .d (n_16099), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[0]));
  CDN_flop \sh_bit_cnt_reg[1] (.clk (clk), .d (n_24624), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[1]));
  CDN_flop \sh_bit_cnt_reg[2] (.clk (clk), .d (n_24590), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[2]));
  CDN_flop \sh_bit_cnt_reg[3] (.clk (clk), .d (n_17057), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_bit_cnt[3]));
  CDN_flop \sh_reg_in_reg[0] (.clk (clk), .d (din), .sena (n_16075),
       .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd (1'b0), .q
       (sh_reg_in[0]));
  CDN_flop \sh_reg_in_reg[1] (.clk (clk), .d (sh_reg_in[0]), .sena
       (n_16075), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (sh_reg_in[1]));
  CDN_flop \sh_reg_in_reg[2] (.clk (clk), .d (sh_reg_in[1]), .sena
       (n_16075), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (sh_reg_in[2]));
  CDN_flop \sh_reg_in_reg[3] (.clk (clk), .d (sh_reg_in[2]), .sena
       (n_16075), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (sh_reg_in[3]));
  CDN_flop \sh_reg_in_reg[4] (.clk (clk), .d (sh_reg_in[3]), .sena
       (n_16075), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (sh_reg_in[4]));
  CDN_flop \sh_reg_in_reg[5] (.clk (clk), .d (sh_reg_in[4]), .sena
       (n_16075), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (sh_reg_in[5]));
  CDN_flop \sh_reg_in_reg[6] (.clk (clk), .d (sh_reg_in[5]), .sena
       (n_16075), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (sh_reg_in[6]));
  CDN_flop \sh_reg_in_reg[7] (.clk (clk), .d (sh_reg_in[6]), .sena
       (n_16075), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (sh_reg_in[7]));
  CDN_flop \sh_reg_in_reg[8] (.clk (clk), .d (sh_reg_in[7]), .sena
       (n_16075), .aclr (1'b0), .apre (1'b0), .srl (n_16074), .srd
       (1'b0), .q (sh_reg_in[8]));
  CDN_flop \sh_reg_out_bit_counter_reg[0] (.clk (clk), .d (n_16107),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[0]));
  CDN_flop \sh_reg_out_bit_counter_reg[1] (.clk (clk), .d (n_24623),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[1]));
  CDN_flop \sh_reg_out_bit_counter_reg[2] (.clk (clk), .d (n_17065),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[2]));
  CDN_flop \sh_reg_out_bit_counter_reg[3] (.clk (clk), .d (n_17064),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[3]));
  CDN_flop \sh_reg_out_bit_counter_reg[4] (.clk (clk), .d (n_17063),
       .sena (1'b1), .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd
       (1'b0), .q (sh_reg_out_bit_counter[4]));
  CDN_flop \sh_reg_out_reg[0] (.clk (clk), .d (n_17080), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[0]));
  CDN_flop \sh_reg_out_reg[1] (.clk (clk), .d (n_17139), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[1]));
  CDN_flop \sh_reg_out_reg[2] (.clk (clk), .d (n_17140), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[2]));
  CDN_flop \sh_reg_out_reg[3] (.clk (clk), .d (n_17141), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[3]));
  CDN_flop \sh_reg_out_reg[4] (.clk (clk), .d (n_17142), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[4]));
  CDN_flop \sh_reg_out_reg[5] (.clk (clk), .d (n_17143), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[5]));
  CDN_flop \sh_reg_out_reg[6] (.clk (clk), .d (n_17144), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[6]));
  CDN_flop \sh_reg_out_reg[7] (.clk (clk), .d (n_17145), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[7]));
  CDN_flop \sh_reg_out_reg[8] (.clk (clk), .d (n_17146), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[8]));
  CDN_flop \sh_reg_out_reg[9] (.clk (clk), .d (n_24625), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[9]));
  CDN_flop \sh_reg_out_reg[10] (.clk (clk), .d (n_17138), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[10]));
  CDN_flop \sh_reg_out_reg[11] (.clk (clk), .d (n_17126), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[11]));
  CDN_flop \sh_reg_out_reg[12] (.clk (clk), .d (n_17130), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[12]));
  CDN_flop \sh_reg_out_reg[13] (.clk (clk), .d (n_17127), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[13]));
  CDN_flop \sh_reg_out_reg[14] (.clk (clk), .d (n_17128), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[14]));
  CDN_flop \sh_reg_out_reg[15] (.clk (clk), .d (n_17129), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[15]));
  CDN_flop \sh_reg_out_reg[16] (.clk (clk), .d (n_17136), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[16]));
  CDN_flop \sh_reg_out_reg[17] (.clk (clk), .d (n_17131), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[17]));
  CDN_flop \sh_reg_out_reg[18] (.clk (clk), .d (n_17132), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[18]));
  CDN_flop \sh_reg_out_reg[19] (.clk (clk), .d (n_24626), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[19]));
  CDN_flop \sh_reg_out_reg[20] (.clk (clk), .d (n_17137), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[20]));
  CDN_flop \sh_reg_out_reg[21] (.clk (clk), .d (n_17147), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[21]));
  CDN_flop \sh_reg_out_reg[22] (.clk (clk), .d (n_24627), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[22]));
  CDN_flop \sh_reg_out_reg[23] (.clk (clk), .d (n_24644), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[23]));
  CDN_flop \sh_reg_out_reg[24] (.clk (clk), .d (n_24609), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[24]));
  CDN_flop \sh_reg_out_reg[25] (.clk (clk), .d (n_24603), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[25]));
  CDN_flop \sh_reg_out_reg[26] (.clk (clk), .d (n_17135), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[26]));
  CDN_flop \sh_reg_out_reg[27] (.clk (clk), .d (n_24604), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[27]));
  CDN_flop \sh_reg_out_reg[28] (.clk (clk), .d (n_17133), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q
       (sh_reg_out[28]));
  CDN_flop \sh_reg_out_reg[29] (.clk (clk), .d (n_17134), .sena (1'b1),
       .aclr (1'b0), .apre (1'b0), .srl (1'b0), .srd (1'b0), .q (dout));
endmodule

`ifdef RC_CDN_GENERIC_GATE
`else
module CDN_flop(clk, d, sena, aclr, apre, srl, srd, q);
  input clk, d, sena, aclr, apre, srl, srd;
  output q;
  wire clk, d, sena, aclr, apre, srl, srd;
  wire q;
  reg  qi;
  assign #1 q = qi;
  always 
    @(posedge clk or posedge apre or posedge aclr) 
      if (aclr) 
        qi <= 0;
      else if (apre) 
          qi <= 1;
        else if (srl) 
            qi <= srd;
          else begin
            if (sena) 
              qi <= d;
          end
  initial 
    qi <= 1'b0;
endmodule
`endif
